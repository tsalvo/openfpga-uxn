-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity dei_0CLK_d0894221 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dei_0CLK_d0894221;
architecture arch of dei_0CLK_d0894221 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal has_written_to_t : unsigned(0 downto 0) := to_unsigned(0, 1);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal device_in_result : device_in_result_t := device_in_result_t_NULL;
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_has_written_to_t : unsigned(0 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_device_in_result : device_in_result_t;
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l401_c6_14c6]
signal BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l411_c7_37df]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l401_c2_82fe]
signal has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l401_c2_82fe]
signal device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : device_in_result_t;

-- result_u8_value_MUX[uxn_opcodes_h_l401_c2_82fe]
signal result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l401_c2_82fe]
signal result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l401_c2_82fe]
signal result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l401_c2_82fe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l401_c2_82fe]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l401_c2_82fe]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l401_c2_82fe]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l401_c2_82fe]
signal t8_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l411_c11_8561]
signal BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l415_c1_06ab]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l411_c7_37df]
signal has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l411_c7_37df]
signal device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_return_output : device_in_result_t;

-- result_u8_value_MUX[uxn_opcodes_h_l411_c7_37df]
signal result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l411_c7_37df]
signal result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l411_c7_37df]
signal result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l411_c7_37df]
signal result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l411_c7_37df]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l411_c7_37df]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l411_c7_37df]
signal t8_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l413_c30_471a]
signal sp_relative_shift_uxn_opcodes_h_l413_c30_471a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l413_c30_471a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l413_c30_471a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l413_c30_471a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l417_c9_b062]
signal BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l417_c9_1e7e]
signal MUX_uxn_opcodes_h_l417_c9_1e7e_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l417_c9_1e7e_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l417_c9_1e7e_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l417_c9_1e7e_return_output : unsigned(7 downto 0);

-- UNARY_OP_NOT[uxn_opcodes_h_l418_c8_8eb4]
signal UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l418_c1_8c9b]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l418_c3_1d50]
signal has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l418_c3_1d50]
signal device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : device_in_result_t;

-- result_u8_value_MUX[uxn_opcodes_h_l418_c3_1d50]
signal result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l418_c3_1d50]
signal result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l418_c3_1d50]
signal result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l418_c3_1d50]
signal result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l418_c3_1d50]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l419_c37_8272]
signal BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_right : unsigned(1 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_return_output : unsigned(7 downto 0);

-- device_in[uxn_opcodes_h_l419_c23_a0ec]
signal device_in_uxn_opcodes_h_l419_c23_a0ec_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_in_uxn_opcodes_h_l419_c23_a0ec_device_address : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l419_c23_a0ec_phase : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l419_c23_a0ec_previous_device_ram_read : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l419_c23_a0ec_return_output : device_in_result_t;

-- UNARY_OP_NOT[uxn_opcodes_h_l422_c9_ef7a]
signal UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l422_c4_f12c]
signal has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l422_c4_f12c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l422_c4_f12c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l422_c4_f12c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l422_c4_f12c]
signal result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_return_output : unsigned(7 downto 0);

function CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6( ref_toks_0 : device_in_result_t;
 ref_toks_1 : unsigned) return device_in_result_t is
 
  variable base : device_in_result_t; 
  variable return_output : device_in_result_t;
begin
      base := ref_toks_0;
      base.is_dei_done := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_ed08( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.device_ram_address := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_device_ram_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6
BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_left,
BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_right,
BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe
has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_cond,
has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe
device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_cond,
device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue,
device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse,
device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe
result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_cond,
result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe
result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe
result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe
result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe
result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe
result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_return_output);

-- t8_MUX_uxn_opcodes_h_l401_c2_82fe
t8_MUX_uxn_opcodes_h_l401_c2_82fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l401_c2_82fe_cond,
t8_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue,
t8_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse,
t8_MUX_uxn_opcodes_h_l401_c2_82fe_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561
BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_left,
BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_right,
BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df
has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_cond,
has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l411_c7_37df
device_in_result_MUX_uxn_opcodes_h_l411_c7_37df : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_cond,
device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iftrue,
device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iffalse,
device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df
result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_cond,
result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df
result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df
result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df
result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df
result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_return_output);

-- t8_MUX_uxn_opcodes_h_l411_c7_37df
t8_MUX_uxn_opcodes_h_l411_c7_37df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l411_c7_37df_cond,
t8_MUX_uxn_opcodes_h_l411_c7_37df_iftrue,
t8_MUX_uxn_opcodes_h_l411_c7_37df_iffalse,
t8_MUX_uxn_opcodes_h_l411_c7_37df_return_output);

-- sp_relative_shift_uxn_opcodes_h_l413_c30_471a
sp_relative_shift_uxn_opcodes_h_l413_c30_471a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l413_c30_471a_ins,
sp_relative_shift_uxn_opcodes_h_l413_c30_471a_x,
sp_relative_shift_uxn_opcodes_h_l413_c30_471a_y,
sp_relative_shift_uxn_opcodes_h_l413_c30_471a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062
BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_left,
BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_right,
BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_return_output);

-- MUX_uxn_opcodes_h_l417_c9_1e7e
MUX_uxn_opcodes_h_l417_c9_1e7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l417_c9_1e7e_cond,
MUX_uxn_opcodes_h_l417_c9_1e7e_iftrue,
MUX_uxn_opcodes_h_l417_c9_1e7e_iffalse,
MUX_uxn_opcodes_h_l417_c9_1e7e_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4
UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_expr,
UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50
has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_cond,
has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50
device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_cond,
device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue,
device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse,
device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50
result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_cond,
result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50
result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50
result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50
result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272
BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272 : entity work.BIN_OP_MINUS_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_left,
BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_right,
BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_return_output);

-- device_in_uxn_opcodes_h_l419_c23_a0ec
device_in_uxn_opcodes_h_l419_c23_a0ec : entity work.device_in_0CLK_85463cfa port map (
clk,
device_in_uxn_opcodes_h_l419_c23_a0ec_CLOCK_ENABLE,
device_in_uxn_opcodes_h_l419_c23_a0ec_device_address,
device_in_uxn_opcodes_h_l419_c23_a0ec_phase,
device_in_uxn_opcodes_h_l419_c23_a0ec_previous_device_ram_read,
device_in_uxn_opcodes_h_l419_c23_a0ec_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a
UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_expr,
UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c
has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_cond,
has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c
result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c
result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c
result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_cond,
result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_device_ram_read,
 -- Registers
 has_written_to_t,
 t8,
 device_in_result,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
 device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
 t8_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_return_output,
 device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_return_output,
 t8_MUX_uxn_opcodes_h_l411_c7_37df_return_output,
 sp_relative_shift_uxn_opcodes_h_l413_c30_471a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_return_output,
 MUX_uxn_opcodes_h_l417_c9_1e7e_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_return_output,
 device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_return_output,
 device_in_uxn_opcodes_h_l419_c23_a0ec_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : device_in_result_t;
 variable VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l401_c2_82fe_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l406_c3_6d35 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_TRUE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l401_c2_82fe_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l416_c3_187e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l418_c8_ba28_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_cond : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_device_address : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_phase : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_return_output : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_return_output : device_in_result_t;
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l420_c32_0c33_return_output : unsigned(7 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l424_c5_d714 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l425_c23_eb92_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l422_l411_l418_l401_DUPLICATE_d72d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_d3f9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_7403_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_5346_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_8ae2_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ed08_uxn_opcodes_h_l395_l434_DUPLICATE_9e30_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_has_written_to_t : unsigned(0 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_device_in_result : device_in_result_t;
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_has_written_to_t := has_written_to_t;
  REG_VAR_t8 := t8;
  REG_VAR_device_in_result := device_in_result;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l406_c3_6d35 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l406_c3_6d35;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l416_c3_187e := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iffalse := VAR_result_sp_relative_shift_uxn_opcodes_h_l416_c3_187e;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_right := to_unsigned(1, 1);
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l424_c5_d714 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l424_c5_d714;
     VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_right := to_unsigned(2, 2);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iffalse := VAR_CLOCK_ENABLE;
     VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iftrue := device_in_result;
     VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse := device_in_result;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_expr := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse := has_written_to_t;
     VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_left := VAR_phase;
     VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_iftrue := VAR_previous_stack_read;
     VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_iftrue := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l417_c9_b062] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_left;
     BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_return_output := BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l411_c11_8561] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_left;
     BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output := BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l422_l411_l418_l401_DUPLICATE_d72d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l422_l411_l418_l401_DUPLICATE_d72d_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l413_c30_471a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l413_c30_471a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_ins;
     sp_relative_shift_uxn_opcodes_h_l413_c30_471a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_x;
     sp_relative_shift_uxn_opcodes_h_l413_c30_471a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_return_output := sp_relative_shift_uxn_opcodes_h_l413_c30_471a_return_output;

     -- result_sp_relative_shift_TRUE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     VAR_result_sp_relative_shift_TRUE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l401_c2_82fe_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d[uxn_opcodes_h_l418_c8_ba28] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l418_c8_ba28_return_output := device_in_result.is_dei_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l401_c6_14c6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_left;
     BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output := BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;

     -- result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l401_c2_82fe_return_output := result.is_device_ram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_7403 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_7403_return_output := result.device_ram_address;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_5346 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_5346_return_output := result.is_opc_done;

     -- UNARY_OP_NOT[uxn_opcodes_h_l422_c9_ef7a] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_return_output := UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_return_output;

     -- CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d[uxn_opcodes_h_l425_c23_eb92] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l425_c23_eb92_return_output := device_in_result.dei_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_d3f9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_d3f9_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_8ae2 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_8ae2_return_output := result.stack_address_sp_offset;

     -- device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l401_c2_82fe_return_output := CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6(
     device_in_result,
     to_unsigned(0, 1));

     -- BIN_OP_MINUS[uxn_opcodes_h_l419_c37_8272] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_left;
     BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_return_output := BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l401_c6_14c6_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l411_c11_8561_return_output;
     VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l417_c9_b062_return_output;
     VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_phase := VAR_BIN_OP_MINUS_uxn_opcodes_h_l419_c37_8272_return_output;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_expr := VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l418_c8_ba28_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_5346_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_5346_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_5346_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_d3f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_d3f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_d3f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_8ae2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_8ae2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l422_l411_l418_DUPLICATE_8ae2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l425_c23_eb92_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_7403_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_7403_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l411_l418_l401_DUPLICATE_7403_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l422_l411_l418_l401_DUPLICATE_d72d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l422_l411_l418_l401_DUPLICATE_d72d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l422_l411_l418_l401_DUPLICATE_d72d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l422_l411_l418_l401_DUPLICATE_d72d_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l422_c9_ef7a_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue := VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l401_c2_82fe_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse := VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l401_c2_82fe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue := VAR_result_sp_relative_shift_TRUE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l401_c2_82fe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l413_c30_471a_return_output;
     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;

     -- MUX[uxn_opcodes_h_l417_c9_1e7e] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l417_c9_1e7e_cond <= VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_cond;
     MUX_uxn_opcodes_h_l417_c9_1e7e_iftrue <= VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_iftrue;
     MUX_uxn_opcodes_h_l417_c9_1e7e_iffalse <= VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_return_output := MUX_uxn_opcodes_h_l417_c9_1e7e_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l422_c4_f12c] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_return_output := has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l422_c4_f12c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l422_c4_f12c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_return_output := result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l422_c4_f12c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_return_output;

     -- UNARY_OP_NOT[uxn_opcodes_h_l418_c8_8eb4] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output := UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l422_c4_f12c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l411_c7_37df] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l411_c7_37df] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l411_c7_37df_return_output;
     VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_device_address := VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_iffalse := VAR_MUX_uxn_opcodes_h_l417_c9_1e7e_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l418_c8_8eb4_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l422_c4_f12c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l422_c4_f12c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l422_c4_f12c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l411_c7_37df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l422_c4_f12c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l422_c4_f12c_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l418_c3_1d50] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l418_c3_1d50] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l418_c3_1d50] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_cond;
     result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_return_output := result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;

     -- t8_MUX[uxn_opcodes_h_l411_c7_37df] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l411_c7_37df_cond <= VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_cond;
     t8_MUX_uxn_opcodes_h_l411_c7_37df_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_iftrue;
     t8_MUX_uxn_opcodes_h_l411_c7_37df_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_return_output := t8_MUX_uxn_opcodes_h_l411_c7_37df_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l415_c1_06ab] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l418_c3_1d50] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l418_c3_1d50] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_return_output := has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;

     -- Submodule level 3
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l415_c1_06ab_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse := VAR_t8_MUX_uxn_opcodes_h_l411_c7_37df_return_output;
     -- has_written_to_t_MUX[uxn_opcodes_h_l411_c7_37df] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_return_output := has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l411_c7_37df] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_cond;
     result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_return_output := result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l411_c7_37df] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_return_output;

     -- t8_MUX[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l401_c2_82fe_cond <= VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_cond;
     t8_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue;
     t8_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_return_output := t8_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l411_c7_37df] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l411_c7_37df] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l418_c1_8c9b] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_return_output;

     -- Submodule level 4
     VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l418_c1_8c9b_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l411_c7_37df_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l411_c7_37df_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l411_c7_37df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l411_c7_37df_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l411_c7_37df_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_cond;
     result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_return_output := result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_return_output := has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;

     -- device_in[uxn_opcodes_h_l419_c23_a0ec] LATENCY=0
     -- Clock enable
     device_in_uxn_opcodes_h_l419_c23_a0ec_CLOCK_ENABLE <= VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_CLOCK_ENABLE;
     -- Inputs
     device_in_uxn_opcodes_h_l419_c23_a0ec_device_address <= VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_device_address;
     device_in_uxn_opcodes_h_l419_c23_a0ec_phase <= VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_phase;
     device_in_uxn_opcodes_h_l419_c23_a0ec_previous_device_ram_read <= VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_previous_device_ram_read;
     -- Outputs
     VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_return_output := device_in_uxn_opcodes_h_l419_c23_a0ec_return_output;

     -- Submodule level 5
     VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue := VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_return_output;
     REG_VAR_has_written_to_t := VAR_has_written_to_t_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;
     -- CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d[uxn_opcodes_h_l420_c32_0c33] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l420_c32_0c33_return_output := VAR_device_in_uxn_opcodes_h_l419_c23_a0ec_return_output.device_ram_address;

     -- device_in_result_MUX[uxn_opcodes_h_l418_c3_1d50] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_cond;
     device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_return_output := device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;

     -- Submodule level 6
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l420_c32_0c33_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l418_c3_1d50] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;

     -- device_in_result_MUX[uxn_opcodes_h_l411_c7_37df] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_cond;
     device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_return_output := device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_return_output;

     -- Submodule level 7
     VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l411_c7_37df_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l418_c3_1d50_return_output;
     -- device_in_result_MUX[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_cond;
     device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_return_output := device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l411_c7_37df] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_return_output;

     -- Submodule level 8
     REG_VAR_device_in_result := VAR_device_in_result_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l411_c7_37df_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l401_c2_82fe] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_ed08_uxn_opcodes_h_l395_l434_DUPLICATE_9e30 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ed08_uxn_opcodes_h_l395_l434_DUPLICATE_9e30_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_ed08(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l401_c2_82fe_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l401_c2_82fe_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ed08_uxn_opcodes_h_l395_l434_DUPLICATE_9e30_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ed08_uxn_opcodes_h_l395_l434_DUPLICATE_9e30_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_has_written_to_t <= REG_VAR_has_written_to_t;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_device_in_result <= REG_VAR_device_in_result;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     has_written_to_t <= REG_COMB_has_written_to_t;
     t8 <= REG_COMB_t8;
     device_in_result <= REG_COMB_device_in_result;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
