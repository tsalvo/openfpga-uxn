-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 42
entity swp_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end swp_0CLK_85d5529e;
architecture arch of swp_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2570_c6_9d5a]
signal BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2570_c2_adaf]
signal t8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2570_c2_adaf]
signal n8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2570_c2_adaf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2570_c2_adaf]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2570_c2_adaf]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2570_c2_adaf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2570_c2_adaf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2570_c2_adaf]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2570_c2_adaf]
signal result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2570_c2_adaf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2570_c2_adaf]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2583_c11_819f]
signal BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2583_c7_96cb]
signal t8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2583_c7_96cb]
signal n8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2583_c7_96cb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2583_c7_96cb]
signal result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2583_c7_96cb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2583_c7_96cb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2583_c7_96cb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2586_c11_727b]
signal BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2586_c7_2e08]
signal t8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2586_c7_2e08]
signal n8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2586_c7_2e08]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2586_c7_2e08]
signal result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2586_c7_2e08]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2586_c7_2e08]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2586_c7_2e08]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2589_c11_5795]
signal BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2589_c7_b9cf]
signal n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2589_c7_b9cf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2589_c7_b9cf]
signal result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2589_c7_b9cf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2589_c7_b9cf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2589_c7_b9cf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2591_c30_0a81]
signal sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2596_c11_3e5e]
signal BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2596_c7_9d57]
signal result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2596_c7_9d57]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2596_c7_9d57]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2596_c7_9d57]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a
BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_left,
BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_right,
BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output);

-- t8_MUX_uxn_opcodes_h_l2570_c2_adaf
t8_MUX_uxn_opcodes_h_l2570_c2_adaf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond,
t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue,
t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse,
t8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

-- n8_MUX_uxn_opcodes_h_l2570_c2_adaf
n8_MUX_uxn_opcodes_h_l2570_c2_adaf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond,
n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue,
n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse,
n8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf
result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf
result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf
result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf
result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf
result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf
result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_cond,
result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf
result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f
BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_left,
BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_right,
BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output);

-- t8_MUX_uxn_opcodes_h_l2583_c7_96cb
t8_MUX_uxn_opcodes_h_l2583_c7_96cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond,
t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue,
t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse,
t8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output);

-- n8_MUX_uxn_opcodes_h_l2583_c7_96cb
n8_MUX_uxn_opcodes_h_l2583_c7_96cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond,
n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue,
n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse,
n8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb
result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb
result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_cond,
result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb
result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb
result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b
BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_left,
BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_right,
BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output);

-- t8_MUX_uxn_opcodes_h_l2586_c7_2e08
t8_MUX_uxn_opcodes_h_l2586_c7_2e08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond,
t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue,
t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse,
t8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output);

-- n8_MUX_uxn_opcodes_h_l2586_c7_2e08
n8_MUX_uxn_opcodes_h_l2586_c7_2e08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond,
n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue,
n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse,
n8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08
result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08
result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_cond,
result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08
result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08
result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795
BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_left,
BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_right,
BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output);

-- n8_MUX_uxn_opcodes_h_l2589_c7_b9cf
n8_MUX_uxn_opcodes_h_l2589_c7_b9cf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond,
n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue,
n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse,
n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf
result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf
result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond,
result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf
result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf
result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81
sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_ins,
sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_x,
sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_y,
sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e
BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_left,
BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_right,
BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57
result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_cond,
result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57
result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57
result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output,
 t8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
 n8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output,
 t8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output,
 n8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output,
 t8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output,
 n8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output,
 n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output,
 sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2575_c3_f0a6 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2580_c3_bc3d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2584_c3_fdec : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2593_c3_533c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2597_c3_8ff6 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2598_c3_a1ea : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2570_DUPLICATE_3ed5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2589_DUPLICATE_a669_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2583_l2596_l2586_DUPLICATE_0f3e_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2583_l2586_l2589_DUPLICATE_e54f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2596_l2586_DUPLICATE_a759_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2603_l2566_DUPLICATE_897c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_right := to_unsigned(4, 3);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2597_c3_8ff6 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2597_c3_8ff6;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2598_c3_a1ea := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2598_c3_a1ea;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2575_c3_f0a6 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2575_c3_f0a6;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2580_c3_bc3d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2580_c3_bc3d;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2593_c3_533c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2593_c3_533c;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2584_c3_fdec := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2584_c3_fdec;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2589_c11_5795] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_left;
     BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output := BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2583_l2586_l2589_DUPLICATE_e54f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2583_l2586_l2589_DUPLICATE_e54f_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2589_DUPLICATE_a669 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2589_DUPLICATE_a669_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2570_DUPLICATE_3ed5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2570_DUPLICATE_3ed5_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2596_c11_3e5e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2583_c11_819f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2591_c30_0a81] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_ins;
     sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_x;
     sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_return_output := sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2570_c6_9d5a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2596_l2586_DUPLICATE_a759 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2596_l2586_DUPLICATE_a759_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2583_l2596_l2586_DUPLICATE_0f3e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2583_l2596_l2586_DUPLICATE_0f3e_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2586_c11_727b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2570_c6_9d5a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2583_c11_819f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2586_c11_727b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2589_c11_5795_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2596_c11_3e5e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2583_l2596_l2586_DUPLICATE_0f3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2583_l2596_l2586_DUPLICATE_0f3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2583_l2596_l2586_DUPLICATE_0f3e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2589_DUPLICATE_a669_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2589_DUPLICATE_a669_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2589_DUPLICATE_a669_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2589_DUPLICATE_a669_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2583_l2586_l2589_DUPLICATE_e54f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2583_l2586_l2589_DUPLICATE_e54f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2583_l2586_l2589_DUPLICATE_e54f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2596_l2586_DUPLICATE_a759_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2596_l2586_DUPLICATE_a759_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2570_DUPLICATE_3ed5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2570_DUPLICATE_3ed5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2570_DUPLICATE_3ed5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2583_l2596_l2586_l2570_DUPLICATE_3ed5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2570_c2_adaf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2591_c30_0a81_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2596_c7_9d57] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output;

     -- n8_MUX[uxn_opcodes_h_l2589_c7_b9cf] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond <= VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond;
     n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue;
     n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output := n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2596_c7_9d57] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2596_c7_9d57] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2596_c7_9d57] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output := result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output;

     -- t8_MUX[uxn_opcodes_h_l2586_c7_2e08] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond <= VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond;
     t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue;
     t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output := t8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2589_c7_b9cf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2596_c7_9d57_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;
     -- t8_MUX[uxn_opcodes_h_l2583_c7_96cb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond <= VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond;
     t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue;
     t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output := t8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2589_c7_b9cf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2589_c7_b9cf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2589_c7_b9cf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output := result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;

     -- n8_MUX[uxn_opcodes_h_l2586_c7_2e08] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond <= VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_cond;
     n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue;
     n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output := n8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2586_c7_2e08] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2589_c7_b9cf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2589_c7_b9cf_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2586_c7_2e08] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2586_c7_2e08] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2586_c7_2e08] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output := result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2583_c7_96cb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;

     -- n8_MUX[uxn_opcodes_h_l2583_c7_96cb] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond <= VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_cond;
     n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue;
     n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output := n8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;

     -- t8_MUX[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond <= VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond;
     t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue;
     t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output := t8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2586_c7_2e08] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2586_c7_2e08_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;
     -- n8_MUX[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond <= VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_cond;
     n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue;
     n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output := n8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2583_c7_96cb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2583_c7_96cb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2583_c7_96cb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output := result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2583_c7_96cb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2583_c7_96cb_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2570_c2_adaf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output := result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2603_l2566_DUPLICATE_897c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2603_l2566_DUPLICATE_897c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2570_c2_adaf_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2603_l2566_DUPLICATE_897c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2603_l2566_DUPLICATE_897c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
