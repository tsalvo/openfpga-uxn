-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 41
entity lit2_0CLK_4351dde2 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lit2_0CLK_4351dde2;
architecture arch of lit2_0CLK_4351dde2 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp8_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp8_high : unsigned(7 downto 0);
signal REG_COMB_tmp8_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l224_c6_27cb]
signal BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l224_c2_6dec]
signal tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l224_c2_6dec]
signal tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l224_c2_6dec]
signal result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l224_c2_6dec]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l224_c2_6dec]
signal result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l224_c2_6dec]
signal result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l224_c2_6dec]
signal result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l224_c2_6dec]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l224_c2_6dec]
signal result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l224_c2_6dec]
signal result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l224_c2_6dec]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l224_c2_6dec]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l237_c11_1e53]
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l237_c7_8aab]
signal tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l237_c7_8aab]
signal tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l237_c7_8aab]
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l237_c7_8aab]
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l237_c7_8aab]
signal result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l237_c7_8aab]
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l237_c7_8aab]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l237_c7_8aab]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l237_c7_8aab]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l239_c22_e995]
signal BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l241_c11_3360]
signal BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l241_c7_63ea]
signal tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l241_c7_63ea]
signal tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l241_c7_63ea]
signal result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l241_c7_63ea]
signal result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l241_c7_63ea]
signal result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l241_c7_63ea]
signal result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l241_c7_63ea]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l241_c7_63ea]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l245_c22_f696]
signal BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_right : unsigned(1 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l249_c11_32fc]
signal BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_return_output : unsigned(0 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l249_c7_5509]
signal tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l249_c7_5509]
signal result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l249_c7_5509]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l249_c7_5509]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l249_c7_5509]
signal result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_1a75( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;
      base.is_pc_updated := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb
BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_left,
BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_right,
BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec
tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec
tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec
result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec
result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec
result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec
result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec
result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec
result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec
result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec
result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53
BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_left,
BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_right,
BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab
tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_cond,
tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab
tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_cond,
tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab
result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond,
result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab
result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab
result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995
BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_left,
BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_right,
BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360
BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_left,
BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_right,
BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea
tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_cond,
tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea
tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_cond,
tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea
result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea
result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea
result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond,
result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea
result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond,
result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea
result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696
BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696 : entity work.BIN_OP_PLUS_uint16_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_left,
BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_right,
BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc
BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_left,
BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_right,
BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509
tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_cond,
tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509
result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_cond,
result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509
result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509
result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_ram_read,
 -- Registers
 tmp8_high,
 tmp8_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l233_c3_231d : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l239_c3_bec3 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l238_c3_dcf7 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l237_c7_8aab_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l245_c3_43dc : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l241_c7_63ea_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l246_c3_b052 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l252_c3_5b46 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_7364_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_9432_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l237_l241_l249_DUPLICATE_6ea7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l237_l241_DUPLICATE_93b1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l237_l249_DUPLICATE_53b8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l257_l219_DUPLICATE_de7e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp8_high : unsigned(7 downto 0);
variable REG_VAR_tmp8_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp8_high := tmp8_high;
  REG_VAR_tmp8_low := tmp8_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l252_c3_5b46 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l252_c3_5b46;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l233_c3_231d := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l233_c3_231d;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_right := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l246_c3_b052 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l246_c3_b052;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_right := to_unsigned(2, 2);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l238_c3_dcf7 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l238_c3_dcf7;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_left := VAR_pc;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_left := VAR_pc;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue := VAR_previous_ram_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iftrue := VAR_previous_ram_read;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue := VAR_previous_ram_read;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iftrue := VAR_previous_ram_read;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse := tmp8_high;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iffalse := tmp8_low;
     -- BIN_OP_PLUS[uxn_opcodes_h_l239_c22_e995] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_left;
     BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_return_output := BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l237_l241_DUPLICATE_93b1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l237_l241_DUPLICATE_93b1_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l237_l241_l249_DUPLICATE_6ea7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l237_l241_l249_DUPLICATE_6ea7_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l224_c6_27cb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_left;
     BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output := BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_7364 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_7364_return_output := result.u8_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l224_c2_6dec_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l237_l249_DUPLICATE_53b8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l237_l249_DUPLICATE_53b8_return_output := result.is_pc_updated;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l237_c7_8aab] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l237_c7_8aab_return_output := result.sp_relative_shift;

     -- result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d[uxn_opcodes_h_l241_c7_63ea] LATENCY=0
     VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l241_c7_63ea_return_output := result.u16_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l224_c2_6dec_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l249_c11_32fc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_left;
     BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_return_output := BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_9432 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_9432_return_output := result.stack_address_sp_offset;

     -- BIN_OP_PLUS[uxn_opcodes_h_l245_c22_f696] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_left;
     BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_return_output := BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l237_c11_1e53] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_left;
     BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output := BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l224_c2_6dec_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l241_c11_3360] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_left;
     BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output := BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l224_c6_27cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_1e53_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_3360_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_32fc_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l239_c3_bec3 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_e995_return_output, 16);
     VAR_result_u16_value_uxn_opcodes_h_l245_c3_43dc := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l245_c22_f696_return_output, 16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l237_l241_l249_DUPLICATE_6ea7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l237_l241_l249_DUPLICATE_6ea7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l237_l241_l249_DUPLICATE_6ea7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l237_l249_DUPLICATE_53b8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l237_l249_DUPLICATE_53b8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l237_l241_DUPLICATE_93b1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l237_l241_DUPLICATE_93b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_9432_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_9432_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_9432_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_7364_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_7364_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l237_l224_l249_DUPLICATE_7364_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l224_c2_6dec_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l224_c2_6dec_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l224_c2_6dec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l237_c7_8aab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse := VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l241_c7_63ea_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue := VAR_result_u16_value_uxn_opcodes_h_l239_c3_bec3;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue := VAR_result_u16_value_uxn_opcodes_h_l245_c3_43dc;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l249_c7_5509] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l249_c7_5509] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l249_c7_5509] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l241_c7_63ea] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_cond;
     tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_return_output := tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l237_c7_8aab] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l249_c7_5509] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_cond;
     result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_return_output := result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l249_c7_5509] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_cond;
     tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_return_output := tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l241_c7_63ea] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l241_c7_63ea] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond;
     result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output := result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_5509_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l249_c7_5509_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l249_c7_5509_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l249_c7_5509_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l249_c7_5509_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l241_c7_63ea] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l237_c7_8aab] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_cond;
     tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_return_output := tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l241_c7_63ea] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l241_c7_63ea] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_cond;
     tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_return_output := tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l241_c7_63ea] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_cond;
     result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output := result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l241_c7_63ea] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l237_c7_8aab] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l237_c7_8aab] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond;
     result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output := result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l241_c7_63ea_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l237_c7_8aab] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_cond;
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output := result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l237_c7_8aab] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_cond;
     tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_return_output := tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l237_c7_8aab] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l237_c7_8aab] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l237_c7_8aab] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;
     REG_VAR_tmp8_high := VAR_tmp8_high_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l237_c7_8aab_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l224_c2_6dec] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_cond;
     result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output := result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;

     -- Submodule level 5
     REG_VAR_tmp8_low := VAR_tmp8_low_MUX_uxn_opcodes_h_l224_c2_6dec_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l257_l219_DUPLICATE_de7e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l257_l219_DUPLICATE_de7e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_1a75(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l224_c2_6dec_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l224_c2_6dec_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l257_l219_DUPLICATE_de7e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l257_l219_DUPLICATE_de7e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp8_high <= REG_VAR_tmp8_high;
REG_COMB_tmp8_low <= REG_VAR_tmp8_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp8_high <= REG_COMB_tmp8_high;
     tmp8_low <= REG_COMB_tmp8_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
