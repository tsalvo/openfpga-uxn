-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity jsr_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr_0CLK_fedec265;
architecture arch of jsr_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l733_c6_ba72]
signal BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l733_c2_e497]
signal result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l733_c2_e497]
signal result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l733_c2_e497]
signal result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l733_c2_e497]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l733_c2_e497]
signal result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l733_c2_e497]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l733_c2_e497]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l733_c2_e497]
signal result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l733_c2_e497]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l733_c2_e497]
signal result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l733_c2_e497]
signal t8_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l746_c11_5a0c]
signal BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l746_c7_eaa8]
signal result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l746_c7_eaa8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l746_c7_eaa8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l746_c7_eaa8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l746_c7_eaa8]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l746_c7_eaa8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l746_c7_eaa8]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l746_c7_eaa8]
signal result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l746_c7_eaa8]
signal t8_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l748_c30_7b8b]
signal sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l750_c11_a034]
signal BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l750_c7_d183]
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l750_c7_d183]
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l750_c7_d183]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l750_c7_d183]
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l750_c7_d183]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l750_c7_d183]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l750_c7_d183]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l750_c7_d183]
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l750_c7_d183]
signal t8_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l758_c11_cb2c]
signal BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l758_c7_5cc1]
signal result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l758_c7_5cc1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l758_c7_5cc1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l758_c7_5cc1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l758_c7_5cc1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l758_c7_5cc1]
signal result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : unsigned(7 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l761_c31_4b53]
signal CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l763_c22_a666]
signal BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_return_output : signed(17 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_a906( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.u8_value := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72
BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_left,
BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_right,
BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497
result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_cond,
result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497
result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497
result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497
result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497
result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497
result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497
result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497
result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_cond,
result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

-- t8_MUX_uxn_opcodes_h_l733_c2_e497
t8_MUX_uxn_opcodes_h_l733_c2_e497 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l733_c2_e497_cond,
t8_MUX_uxn_opcodes_h_l733_c2_e497_iftrue,
t8_MUX_uxn_opcodes_h_l733_c2_e497_iffalse,
t8_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c
BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_left,
BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_right,
BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8
result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond,
result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8
result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8
result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8
result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8
result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8
result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond,
result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output);

-- t8_MUX_uxn_opcodes_h_l746_c7_eaa8
t8_MUX_uxn_opcodes_h_l746_c7_eaa8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l746_c7_eaa8_cond,
t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue,
t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse,
t8_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output);

-- sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b
sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_ins,
sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_x,
sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_y,
sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034
BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_left,
BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_right,
BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183
result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_cond,
result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183
result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_cond,
result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output);

-- t8_MUX_uxn_opcodes_h_l750_c7_d183
t8_MUX_uxn_opcodes_h_l750_c7_d183 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l750_c7_d183_cond,
t8_MUX_uxn_opcodes_h_l750_c7_d183_iftrue,
t8_MUX_uxn_opcodes_h_l750_c7_d183_iffalse,
t8_MUX_uxn_opcodes_h_l750_c7_d183_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c
BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_left,
BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_right,
BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1
result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond,
result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1
result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1
result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1
result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1
result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond,
result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output);

-- CONST_SR_8_uxn_opcodes_h_l761_c31_4b53
CONST_SR_8_uxn_opcodes_h_l761_c31_4b53 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_x,
CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666
BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_left,
BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_right,
BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
 t8_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output,
 t8_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output,
 sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output,
 t8_MUX_uxn_opcodes_h_l750_c7_d183_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output,
 CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l743_c3_e565 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l738_c3_6040 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l747_c3_25bf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l755_c3_f2bb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l753_c3_5aca : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l756_c21_64ec_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l763_c3_a4a6 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_b5bf : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l758_c7_5cc1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l760_c3_2305 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l758_c7_5cc1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l761_c21_92a2_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l763_c27_0f40_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_return_output : signed(17 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_9178_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_f7c1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_535c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_df5f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_6b09_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_5f6e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l729_l767_DUPLICATE_ce75_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l760_c3_2305 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l760_c3_2305;
     VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l747_c3_25bf := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l747_c3_25bf;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l738_c3_6040 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l738_c3_6040;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l743_c3_e565 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l743_c3_e565;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_right := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l755_c3_f2bb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l755_c3_f2bb;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_b5bf := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_b5bf;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l753_c3_5aca := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l753_c3_5aca;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l748_c30_7b8b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_ins;
     sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_x;
     sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_return_output := sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l733_c2_e497_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l750_c11_a034] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_left;
     BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output := BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l758_c11_cb2c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_left;
     BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output := BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l746_c11_5a0c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_left;
     BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output := BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_f7c1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_f7c1_return_output := result.u8_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l758_c7_5cc1] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l758_c7_5cc1_return_output := result.stack_address_sp_offset;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l756_c21_64ec] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l756_c21_64ec_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_9178 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_9178_return_output := result.u16_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l733_c2_e497_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_6b09 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_6b09_return_output := result.is_stack_index_flipped;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l758_c7_5cc1] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l758_c7_5cc1_return_output := result.sp_relative_shift;

     -- CONST_SR_8[uxn_opcodes_h_l761_c31_4b53] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_x <= VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_return_output := CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_535c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_535c_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_5f6e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_5f6e_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_df5f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_df5f_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l733_c6_ba72] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_left;
     BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output := BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l763_c27_0f40] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l763_c27_0f40_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l733_c6_ba72_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l746_c11_5a0c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l750_c11_a034_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l758_c11_cb2c_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l763_c27_0f40_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l756_c21_64ec_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_9178_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_9178_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_9178_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l750_l733_l758_l746_DUPLICATE_9178_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_535c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_535c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_535c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_5f6e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_5f6e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l750_l758_l746_DUPLICATE_5f6e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_6b09_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_6b09_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_df5f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l750_l746_DUPLICATE_df5f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_f7c1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_f7c1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l733_l758_l746_DUPLICATE_f7c1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l733_c2_e497_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l733_c2_e497_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l758_c7_5cc1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l758_c7_5cc1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l748_c30_7b8b_return_output;
     -- BIN_OP_PLUS[uxn_opcodes_h_l763_c22_a666] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_left;
     BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_return_output := BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_return_output;

     -- t8_MUX[uxn_opcodes_h_l750_c7_d183] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l750_c7_d183_cond <= VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_cond;
     t8_MUX_uxn_opcodes_h_l750_c7_d183_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_iftrue;
     t8_MUX_uxn_opcodes_h_l750_c7_d183_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_return_output := t8_MUX_uxn_opcodes_h_l750_c7_d183_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l750_c7_d183] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l758_c7_5cc1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l758_c7_5cc1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l750_c7_d183] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l758_c7_5cc1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l758_c7_5cc1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l761_c21_92a2] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l761_c21_92a2_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l761_c31_4b53_return_output);

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l763_c3_a4a6 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l763_c22_a666_return_output)),16);
     VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l761_c21_92a2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l750_c7_d183_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l750_c7_d183_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l750_c7_d183_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue := VAR_result_u16_value_uxn_opcodes_h_l763_c3_a4a6;
     -- result_u8_value_MUX[uxn_opcodes_h_l758_c7_5cc1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output := result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l758_c7_5cc1] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_cond;
     result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output := result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;

     -- t8_MUX[uxn_opcodes_h_l746_c7_eaa8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l746_c7_eaa8_cond <= VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_cond;
     t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue;
     t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output := t8_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l746_c7_eaa8] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l750_c7_d183] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l746_c7_eaa8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l750_c7_d183] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l750_c7_d183] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l750_c7_d183] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l750_c7_d183_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l750_c7_d183_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l750_c7_d183_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l750_c7_d183_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l758_c7_5cc1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_iffalse := VAR_t8_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l746_c7_eaa8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l746_c7_eaa8] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l746_c7_eaa8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;

     -- t8_MUX[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l733_c2_e497_cond <= VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_cond;
     t8_MUX_uxn_opcodes_h_l733_c2_e497_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_iftrue;
     t8_MUX_uxn_opcodes_h_l733_c2_e497_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_return_output := t8_MUX_uxn_opcodes_h_l733_c2_e497_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l750_c7_d183] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_cond;
     result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output := result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l750_c7_d183] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_cond;
     result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output := result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l746_c7_eaa8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l750_c7_d183_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l733_c2_e497_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l746_c7_eaa8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output := result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l746_c7_eaa8] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_cond;
     result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output := result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_return_output;

     -- Submodule level 5
     VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l746_c7_eaa8_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_cond;
     result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output := result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l733_c2_e497] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_cond;
     result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output := result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l729_l767_DUPLICATE_ce75 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l729_l767_DUPLICATE_ce75_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a906(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l733_c2_e497_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l733_c2_e497_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l729_l767_DUPLICATE_ce75_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a906_uxn_opcodes_h_l729_l767_DUPLICATE_ce75_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
