-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 56
entity swp_0CLK_bf6dd460 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end swp_0CLK_bf6dd460;
architecture arch of swp_0CLK_bf6dd460 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2710_c6_5d34]
signal BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2710_c1_26ef]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2710_c2_a99e]
signal n8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2710_c2_a99e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2710_c2_a99e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2710_c2_a99e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2710_c2_a99e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2710_c2_a99e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2710_c2_a99e]
signal result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2710_c2_a99e]
signal t8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2711_c3_6011[uxn_opcodes_h_l2711_c3_6011]
signal printf_uxn_opcodes_h_l2711_c3_6011_uxn_opcodes_h_l2711_c3_6011_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2715_c11_75a5]
signal BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2715_c7_fdc1]
signal n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2715_c7_fdc1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2715_c7_fdc1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2715_c7_fdc1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2715_c7_fdc1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2715_c7_fdc1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2715_c7_fdc1]
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2715_c7_fdc1]
signal t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2718_c11_8f59]
signal BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2718_c7_e42e]
signal n8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2718_c7_e42e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2718_c7_e42e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2718_c7_e42e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2718_c7_e42e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2718_c7_e42e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2718_c7_e42e]
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2718_c7_e42e]
signal t8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2722_c11_2b5a]
signal BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2722_c7_b191]
signal n8_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2722_c7_b191]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2722_c7_b191]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2722_c7_b191]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2722_c7_b191]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2722_c7_b191]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2722_c7_b191]
signal result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2725_c11_c86c]
signal BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2725_c7_8e8a]
signal n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2725_c7_8e8a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2725_c7_8e8a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2725_c7_8e8a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2725_c7_8e8a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2725_c7_8e8a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2725_c7_8e8a]
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2728_c30_f76f]
signal sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2733_c11_22b0]
signal BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2733_c7_da08]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2733_c7_da08]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2733_c7_da08]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2733_c7_da08]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2733_c7_da08]
signal result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2738_c11_c963]
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2738_c7_a137]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2738_c7_a137]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8cda( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34
BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_left,
BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_right,
BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_return_output);

-- n8_MUX_uxn_opcodes_h_l2710_c2_a99e
n8_MUX_uxn_opcodes_h_l2710_c2_a99e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond,
n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue,
n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse,
n8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e
result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e
result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e
result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e
result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output);

-- t8_MUX_uxn_opcodes_h_l2710_c2_a99e
t8_MUX_uxn_opcodes_h_l2710_c2_a99e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond,
t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue,
t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse,
t8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output);

-- printf_uxn_opcodes_h_l2711_c3_6011_uxn_opcodes_h_l2711_c3_6011
printf_uxn_opcodes_h_l2711_c3_6011_uxn_opcodes_h_l2711_c3_6011 : entity work.printf_uxn_opcodes_h_l2711_c3_6011_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2711_c3_6011_uxn_opcodes_h_l2711_c3_6011_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5
BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_left,
BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_right,
BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output);

-- n8_MUX_uxn_opcodes_h_l2715_c7_fdc1
n8_MUX_uxn_opcodes_h_l2715_c7_fdc1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond,
n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue,
n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse,
n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1
result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output);

-- t8_MUX_uxn_opcodes_h_l2715_c7_fdc1
t8_MUX_uxn_opcodes_h_l2715_c7_fdc1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond,
t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue,
t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse,
t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_left,
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_right,
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output);

-- n8_MUX_uxn_opcodes_h_l2718_c7_e42e
n8_MUX_uxn_opcodes_h_l2718_c7_e42e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond,
n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue,
n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse,
n8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output);

-- t8_MUX_uxn_opcodes_h_l2718_c7_e42e
t8_MUX_uxn_opcodes_h_l2718_c7_e42e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond,
t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue,
t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse,
t8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a
BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_left,
BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_right,
BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output);

-- n8_MUX_uxn_opcodes_h_l2722_c7_b191
n8_MUX_uxn_opcodes_h_l2722_c7_b191 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2722_c7_b191_cond,
n8_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue,
n8_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse,
n8_MUX_uxn_opcodes_h_l2722_c7_b191_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191
result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191
result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191
result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191
result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191
result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_cond,
result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_left,
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_right,
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output);

-- n8_MUX_uxn_opcodes_h_l2725_c7_8e8a
n8_MUX_uxn_opcodes_h_l2725_c7_8e8a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond,
n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue,
n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse,
n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f
sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_ins,
sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_x,
sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_y,
sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0
BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_left,
BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_right,
BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08
result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08
result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08
result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08
result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_cond,
result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_left,
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_right,
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_return_output,
 n8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
 t8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output,
 n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output,
 t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output,
 n8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output,
 t8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output,
 n8_MUX_uxn_opcodes_h_l2722_c7_b191_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output,
 n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output,
 sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2712_c3_edb3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2711_c3_6011_uxn_opcodes_h_l2711_c3_6011_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2716_c3_e7a8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2720_c3_69db : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2723_c3_4c63 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2730_c3_6972 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2735_c3_86f8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2733_c7_da08_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2715_l2710_l2725_l2722_l2718_DUPLICATE_7176_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_7167_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2715_l2710_l2738_l2733_l2722_l2718_DUPLICATE_61f8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_0a63_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2715_l2738_l2733_l2725_l2722_l2718_DUPLICATE_6151_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2743_l2706_DUPLICATE_0d26_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2730_c3_6972 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2730_c3_6972;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2735_c3_86f8 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2735_c3_86f8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_right := to_unsigned(3, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2723_c3_4c63 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2723_c3_4c63;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_right := to_unsigned(6, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2720_c3_69db := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2720_c3_69db;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2712_c3_edb3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2712_c3_edb3;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2716_c3_e7a8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2716_c3_e7a8;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2722_c11_2b5a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2728_c30_f76f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_ins;
     sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_x;
     sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_return_output := sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_7167 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_7167_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2733_c11_22b0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2733_c7_da08] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2733_c7_da08_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2715_l2738_l2733_l2725_l2722_l2718_DUPLICATE_6151 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2715_l2738_l2733_l2725_l2722_l2718_DUPLICATE_6151_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2715_l2710_l2738_l2733_l2722_l2718_DUPLICATE_61f8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2715_l2710_l2738_l2733_l2722_l2718_DUPLICATE_61f8_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2718_c11_8f59] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_left;
     BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output := BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2710_c6_5d34] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_left;
     BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output := BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2725_c11_c86c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2715_c11_75a5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2738_c11_c963] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_left;
     BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_return_output := BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_0a63 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_0a63_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2715_l2710_l2725_l2722_l2718_DUPLICATE_7176 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2715_l2710_l2725_l2722_l2718_DUPLICATE_7176_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_5d34_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_75a5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_8f59_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_2b5a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_c86c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_22b0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_c963_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2715_l2710_l2725_l2722_l2718_DUPLICATE_7176_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2715_l2710_l2725_l2722_l2718_DUPLICATE_7176_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2715_l2710_l2725_l2722_l2718_DUPLICATE_7176_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2715_l2710_l2725_l2722_l2718_DUPLICATE_7176_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2715_l2710_l2725_l2722_l2718_DUPLICATE_7176_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2715_l2738_l2733_l2725_l2722_l2718_DUPLICATE_6151_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2715_l2738_l2733_l2725_l2722_l2718_DUPLICATE_6151_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2715_l2738_l2733_l2725_l2722_l2718_DUPLICATE_6151_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2715_l2738_l2733_l2725_l2722_l2718_DUPLICATE_6151_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2715_l2738_l2733_l2725_l2722_l2718_DUPLICATE_6151_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2715_l2738_l2733_l2725_l2722_l2718_DUPLICATE_6151_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_7167_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_7167_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_7167_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_7167_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_7167_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2715_l2710_l2738_l2733_l2722_l2718_DUPLICATE_61f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2715_l2710_l2738_l2733_l2722_l2718_DUPLICATE_61f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2715_l2710_l2738_l2733_l2722_l2718_DUPLICATE_61f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2715_l2710_l2738_l2733_l2722_l2718_DUPLICATE_61f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2715_l2710_l2738_l2733_l2722_l2718_DUPLICATE_61f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2715_l2710_l2738_l2733_l2722_l2718_DUPLICATE_61f8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_0a63_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_0a63_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_0a63_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_0a63_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2715_l2710_l2733_l2722_l2718_DUPLICATE_0a63_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2733_c7_da08_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_f76f_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2733_c7_da08] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2710_c1_26ef] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2733_c7_da08] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_return_output := result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_return_output;

     -- t8_MUX[uxn_opcodes_h_l2718_c7_e42e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond;
     t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue;
     t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output := t8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2725_c7_8e8a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2733_c7_da08] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2738_c7_a137] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2738_c7_a137] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_return_output;

     -- n8_MUX[uxn_opcodes_h_l2725_c7_8e8a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond;
     n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue;
     n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output := n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2711_c3_6011_uxn_opcodes_h_l2711_c3_6011_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_26ef_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_a137_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_da08_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_a137_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_da08_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_da08_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;
     -- t8_MUX[uxn_opcodes_h_l2715_c7_fdc1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond <= VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond;
     t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue;
     t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output := t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2725_c7_8e8a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2733_c7_da08] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_return_output;

     -- printf_uxn_opcodes_h_l2711_c3_6011[uxn_opcodes_h_l2711_c3_6011] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2711_c3_6011_uxn_opcodes_h_l2711_c3_6011_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2711_c3_6011_uxn_opcodes_h_l2711_c3_6011_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2733_c7_da08] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_return_output;

     -- n8_MUX[uxn_opcodes_h_l2722_c7_b191] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2722_c7_b191_cond <= VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_cond;
     n8_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue;
     n8_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_return_output := n8_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2725_c7_8e8a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2722_c7_b191] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2725_c7_8e8a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_da08_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_da08_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;
     -- t8_MUX[uxn_opcodes_h_l2710_c2_a99e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond;
     t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue;
     t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output := t8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2725_c7_8e8a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2722_c7_b191] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2722_c7_b191] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2718_c7_e42e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2722_c7_b191] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_return_output := result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2725_c7_8e8a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;

     -- n8_MUX[uxn_opcodes_h_l2718_c7_e42e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond <= VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_cond;
     n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue;
     n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output := n8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_8e8a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2722_c7_b191] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;

     -- n8_MUX[uxn_opcodes_h_l2715_c7_fdc1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond <= VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond;
     n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue;
     n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output := n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2718_c7_e42e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2718_c7_e42e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2718_c7_e42e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2722_c7_b191] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2715_c7_fdc1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_b191_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2710_c2_a99e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2718_c7_e42e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2710_c2_a99e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond <= VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_cond;
     n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue;
     n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output := n8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2715_c7_fdc1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2715_c7_fdc1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2715_c7_fdc1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2718_c7_e42e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_e42e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2710_c2_a99e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2715_c7_fdc1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2715_c7_fdc1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2710_c2_a99e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2710_c2_a99e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_fdc1_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2710_c2_a99e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2710_c2_a99e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2743_l2706_DUPLICATE_0d26 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2743_l2706_DUPLICATE_0d26_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8cda(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_a99e_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2743_l2706_DUPLICATE_0d26_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l2743_l2706_DUPLICATE_0d26_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
