-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity jsr_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr_0CLK_f62d646e;
architecture arch of jsr_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l700_c6_10a1]
signal BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l700_c2_4163]
signal result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l700_c2_4163]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l700_c2_4163]
signal result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l700_c2_4163]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l700_c2_4163]
signal result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l700_c2_4163]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l700_c2_4163]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l700_c2_4163]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l700_c2_4163]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l700_c2_4163]
signal t8_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l707_c11_dfab]
signal BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l707_c7_96a4]
signal result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l707_c7_96a4]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l707_c7_96a4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l707_c7_96a4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l707_c7_96a4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l707_c7_96a4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l707_c7_96a4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l707_c7_96a4]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l707_c7_96a4]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l707_c7_96a4]
signal t8_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l710_c30_9298]
signal sp_relative_shift_uxn_opcodes_h_l710_c30_9298_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l710_c30_9298_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l710_c30_9298_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l710_c30_9298_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l712_c11_cd25]
signal BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l712_c7_2f5f]
signal result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l712_c7_2f5f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l712_c7_2f5f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l712_c7_2f5f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l712_c7_2f5f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l712_c7_2f5f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l712_c7_2f5f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l712_c7_2f5f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l712_c7_2f5f]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l712_c7_2f5f]
signal t8_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l721_c11_6949]
signal BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l721_c7_2580]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l721_c7_2580]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l721_c7_2580]
signal result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(15 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l721_c7_2580]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l721_c7_2580]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l721_c7_2580]
signal result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l721_c7_2580]
signal result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l726_c22_050e]
signal BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l728_c11_ae78]
signal BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l728_c7_982e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l728_c7_982e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l728_c7_982e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_4b08( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_sp_shift := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_stack_operation_16bit := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1
BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_left,
BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_right,
BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163
result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_cond,
result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163
result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163
result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163
result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163
result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163
result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_return_output);

-- t8_MUX_uxn_opcodes_h_l700_c2_4163
t8_MUX_uxn_opcodes_h_l700_c2_4163 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l700_c2_4163_cond,
t8_MUX_uxn_opcodes_h_l700_c2_4163_iftrue,
t8_MUX_uxn_opcodes_h_l700_c2_4163_iffalse,
t8_MUX_uxn_opcodes_h_l700_c2_4163_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab
BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_left,
BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_right,
BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4
result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_cond,
result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4
result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4
result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4
result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4
result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4
result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_return_output);

-- t8_MUX_uxn_opcodes_h_l707_c7_96a4
t8_MUX_uxn_opcodes_h_l707_c7_96a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l707_c7_96a4_cond,
t8_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue,
t8_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse,
t8_MUX_uxn_opcodes_h_l707_c7_96a4_return_output);

-- sp_relative_shift_uxn_opcodes_h_l710_c30_9298
sp_relative_shift_uxn_opcodes_h_l710_c30_9298 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l710_c30_9298_ins,
sp_relative_shift_uxn_opcodes_h_l710_c30_9298_x,
sp_relative_shift_uxn_opcodes_h_l710_c30_9298_y,
sp_relative_shift_uxn_opcodes_h_l710_c30_9298_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25
BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_left,
BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_right,
BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f
result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_cond,
result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f
result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f
result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f
result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f
result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f
result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output);

-- t8_MUX_uxn_opcodes_h_l712_c7_2f5f
t8_MUX_uxn_opcodes_h_l712_c7_2f5f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l712_c7_2f5f_cond,
t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue,
t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse,
t8_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949
BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_left,
BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_right,
BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580
result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580
result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_cond,
result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580
result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580
result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580
result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e
BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_left,
BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_right,
BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78
BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_left,
BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_right,
BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e
result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e
result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
 t8_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_return_output,
 t8_MUX_uxn_opcodes_h_l707_c7_96a4_return_output,
 sp_relative_shift_uxn_opcodes_h_l710_c30_9298_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output,
 t8_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l704_c3_05c7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l708_c3_79f9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l715_c3_0f55 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l717_c3_18d8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l712_c7_2f5f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l726_c3_fa86 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l726_c27_b29c_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_f31e_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l707_l728_l712_l700_DUPLICATE_64e4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l712_l700_DUPLICATE_fb51_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_ee04_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l700_l721_DUPLICATE_e013_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l707_l728_l700_l721_DUPLICATE_490f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_af4c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l707_l728_l712_l721_DUPLICATE_9593_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4b08_uxn_opcodes_h_l696_l734_DUPLICATE_fac9_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l715_c3_0f55 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l715_c3_0f55;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l717_c3_18d8 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l717_c3_18d8;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l708_c3_79f9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l708_c3_79f9;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l704_c3_05c7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l704_c3_05c7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l710_c30_9298] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l710_c30_9298_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_ins;
     sp_relative_shift_uxn_opcodes_h_l710_c30_9298_x <= VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_x;
     sp_relative_shift_uxn_opcodes_h_l710_c30_9298_y <= VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_return_output := sp_relative_shift_uxn_opcodes_h_l710_c30_9298_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l712_c7_2f5f] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l712_c7_2f5f_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_ee04 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_ee04_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l700_l721_DUPLICATE_e013 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l700_l721_DUPLICATE_e013_return_output := result.is_sp_shift;

     -- CAST_TO_int8_t[uxn_opcodes_h_l726_c27_b29c] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l726_c27_b29c_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- BIN_OP_EQ[uxn_opcodes_h_l728_c11_ae78] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_left;
     BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_return_output := BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l707_l728_l712_l700_DUPLICATE_64e4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l707_l728_l712_l700_DUPLICATE_64e4_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l700_c6_10a1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_left;
     BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output := BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l712_c11_cd25] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_left;
     BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output := BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l721_c11_6949] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_left;
     BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output := BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l712_l700_DUPLICATE_fb51 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l712_l700_DUPLICATE_fb51_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_f31e LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_f31e_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l707_l728_l712_l721_DUPLICATE_9593 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l707_l728_l712_l721_DUPLICATE_9593_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l707_l728_l700_l721_DUPLICATE_490f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l707_l728_l700_l721_DUPLICATE_490f_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l707_c11_dfab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_left;
     BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output := BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_af4c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_af4c_return_output := result.is_stack_operation_16bit;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l700_c6_10a1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c11_dfab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c11_cd25_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l721_c11_6949_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l728_c11_ae78_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l726_c27_b29c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l712_l700_DUPLICATE_fb51_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l712_l700_DUPLICATE_fb51_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_f31e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_f31e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_f31e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l707_l728_l712_l721_DUPLICATE_9593_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l707_l728_l712_l721_DUPLICATE_9593_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l707_l728_l712_l721_DUPLICATE_9593_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l707_l728_l712_l721_DUPLICATE_9593_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l707_l728_l712_l700_DUPLICATE_64e4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l707_l728_l712_l700_DUPLICATE_64e4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l707_l728_l712_l700_DUPLICATE_64e4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l707_l728_l712_l700_DUPLICATE_64e4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l700_l721_DUPLICATE_e013_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l700_l721_DUPLICATE_e013_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l700_l721_DUPLICATE_e013_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l707_l728_l700_l721_DUPLICATE_490f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l707_l728_l700_l721_DUPLICATE_490f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l707_l728_l700_l721_DUPLICATE_490f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l707_l728_l700_l721_DUPLICATE_490f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_af4c_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_af4c_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_af4c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_ee04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_ee04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l707_l700_l721_DUPLICATE_ee04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l712_c7_2f5f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l710_c30_9298_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l712_c7_2f5f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l712_c7_2f5f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l728_c7_982e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l728_c7_982e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l721_c7_2580] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l726_c22_050e] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_left;
     BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_return_output := BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l721_c7_2580] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_return_output;

     -- t8_MUX[uxn_opcodes_h_l712_c7_2f5f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l712_c7_2f5f_cond <= VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_cond;
     t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue;
     t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output := t8_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l721_c7_2580] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l728_c7_982e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l726_c3_fa86 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l726_c22_050e_return_output)),16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l728_c7_982e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l728_c7_982e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l721_c7_2580_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l728_c7_982e_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l721_c7_2580_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l721_c7_2580_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iftrue := VAR_result_u16_value_uxn_opcodes_h_l726_c3_fa86;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l707_c7_96a4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l721_c7_2580] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l721_c7_2580] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_cond;
     result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_return_output := result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l721_c7_2580] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l712_c7_2f5f] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l712_c7_2f5f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;

     -- t8_MUX[uxn_opcodes_h_l707_c7_96a4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l707_c7_96a4_cond <= VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_cond;
     t8_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue;
     t8_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_return_output := t8_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l712_c7_2f5f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l721_c7_2580] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l707_c7_96a4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l721_c7_2580_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l721_c7_2580_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l721_c7_2580_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l721_c7_2580_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_iffalse := VAR_t8_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l712_c7_2f5f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l707_c7_96a4] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l707_c7_96a4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l700_c2_4163] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l707_c7_96a4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l700_c2_4163] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l712_c7_2f5f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output := result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l712_c7_2f5f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l712_c7_2f5f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;

     -- t8_MUX[uxn_opcodes_h_l700_c2_4163] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l700_c2_4163_cond <= VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_cond;
     t8_MUX_uxn_opcodes_h_l700_c2_4163_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_iftrue;
     t8_MUX_uxn_opcodes_h_l700_c2_4163_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_return_output := t8_MUX_uxn_opcodes_h_l700_c2_4163_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c7_2f5f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l700_c2_4163_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l707_c7_96a4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l700_c2_4163] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l700_c2_4163] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l700_c2_4163] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l707_c7_96a4] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_cond;
     result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_return_output := result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l707_c7_96a4] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l707_c7_96a4] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l707_c7_96a4_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l700_c2_4163] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l700_c2_4163] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l700_c2_4163] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_cond;
     result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_return_output := result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l700_c2_4163] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4b08_uxn_opcodes_h_l696_l734_DUPLICATE_fac9 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4b08_uxn_opcodes_h_l696_l734_DUPLICATE_fac9_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4b08(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l700_c2_4163_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l700_c2_4163_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4b08_uxn_opcodes_h_l696_l734_DUPLICATE_fac9_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4b08_uxn_opcodes_h_l696_l734_DUPLICATE_fac9_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
