-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity equ_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_226c8821;
architecture arch of equ_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1163_c6_39db]
signal BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1163_c2_1dfb]
signal n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1163_c2_1dfb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1163_c2_1dfb]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1163_c2_1dfb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1163_c2_1dfb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1163_c2_1dfb]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1163_c2_1dfb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1163_c2_1dfb]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1163_c2_1dfb]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1163_c2_1dfb]
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1163_c2_1dfb]
signal t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1176_c11_df2f]
signal BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1176_c7_04de]
signal n8_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1176_c7_04de]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1176_c7_04de]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1176_c7_04de]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1176_c7_04de]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1176_c7_04de]
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1176_c7_04de]
signal t8_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1179_c11_3e50]
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1179_c7_4023]
signal n8_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1179_c7_4023]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1179_c7_4023]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1179_c7_4023]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1179_c7_4023]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1179_c7_4023]
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1179_c7_4023]
signal t8_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1182_c11_f448]
signal BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1182_c7_80b2]
signal n8_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1182_c7_80b2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1182_c7_80b2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1182_c7_80b2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1182_c7_80b2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1182_c7_80b2]
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1184_c30_6ea6]
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1187_c21_ac77]
signal BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1187_c21_9865]
signal MUX_uxn_opcodes_h_l1187_c21_9865_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1187_c21_9865_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1187_c21_9865_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1187_c21_9865_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_04b4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_left,
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_right,
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output);

-- n8_MUX_uxn_opcodes_h_l1163_c2_1dfb
n8_MUX_uxn_opcodes_h_l1163_c2_1dfb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond,
n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue,
n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse,
n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond,
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

-- t8_MUX_uxn_opcodes_h_l1163_c2_1dfb
t8_MUX_uxn_opcodes_h_l1163_c2_1dfb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond,
t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue,
t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse,
t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_left,
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_right,
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output);

-- n8_MUX_uxn_opcodes_h_l1176_c7_04de
n8_MUX_uxn_opcodes_h_l1176_c7_04de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1176_c7_04de_cond,
n8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue,
n8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse,
n8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_cond,
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_return_output);

-- t8_MUX_uxn_opcodes_h_l1176_c7_04de
t8_MUX_uxn_opcodes_h_l1176_c7_04de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1176_c7_04de_cond,
t8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue,
t8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse,
t8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_left,
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_right,
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output);

-- n8_MUX_uxn_opcodes_h_l1179_c7_4023
n8_MUX_uxn_opcodes_h_l1179_c7_4023 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1179_c7_4023_cond,
n8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue,
n8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse,
n8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_cond,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_return_output);

-- t8_MUX_uxn_opcodes_h_l1179_c7_4023
t8_MUX_uxn_opcodes_h_l1179_c7_4023 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1179_c7_4023_cond,
t8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue,
t8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse,
t8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_left,
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_right,
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output);

-- n8_MUX_uxn_opcodes_h_l1182_c7_80b2
n8_MUX_uxn_opcodes_h_l1182_c7_80b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1182_c7_80b2_cond,
n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue,
n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse,
n8_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6
sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_ins,
sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_x,
sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_y,
sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_left,
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_right,
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_return_output);

-- MUX_uxn_opcodes_h_l1187_c21_9865
MUX_uxn_opcodes_h_l1187_c21_9865 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1187_c21_9865_cond,
MUX_uxn_opcodes_h_l1187_c21_9865_iftrue,
MUX_uxn_opcodes_h_l1187_c21_9865_iffalse,
MUX_uxn_opcodes_h_l1187_c21_9865_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output,
 n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
 t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output,
 n8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_return_output,
 t8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output,
 n8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_return_output,
 t8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output,
 n8_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output,
 sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_return_output,
 MUX_uxn_opcodes_h_l1187_c21_9865_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1173_c3_243e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1168_c3_7f4e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1177_c3_e03f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_a798 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_9865_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_9865_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_9865_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_9865_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_8378_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_6a5b_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_536c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_121e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1182_l1179_DUPLICATE_afe6_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1191_l1159_DUPLICATE_19d0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_a798 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_a798;
     VAR_MUX_uxn_opcodes_h_l1187_c21_9865_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1168_c3_7f4e := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1168_c3_7f4e;
     VAR_MUX_uxn_opcodes_h_l1187_c21_9865_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1173_c3_243e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1173_c3_243e;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1177_c3_e03f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1177_c3_e03f;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_6a5b LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_6a5b_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1182_c11_f448] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_left;
     BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output := BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_536c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_536c_return_output := result.is_opc_done;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1179_c11_3e50] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_left;
     BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output := BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output := result.is_ram_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_121e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_121e_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l1184_c30_6ea6] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_ins;
     sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_x;
     sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_return_output := sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1182_l1179_DUPLICATE_afe6 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1182_l1179_DUPLICATE_afe6_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1163_c6_39db] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_left;
     BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output := BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1176_c11_df2f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_8378 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_8378_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1187_c21_ac77] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_left;
     BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_return_output := BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output := result.is_stack_index_flipped;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_39db_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_df2f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_3e50_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_f448_return_output;
     VAR_MUX_uxn_opcodes_h_l1187_c21_9865_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_ac77_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_6a5b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_6a5b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_6a5b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_536c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_536c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_536c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_121e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_121e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1182_l1176_l1179_DUPLICATE_121e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1182_l1179_DUPLICATE_afe6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1182_l1179_DUPLICATE_afe6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_8378_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_8378_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_8378_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1163_l1182_l1176_l1179_DUPLICATE_8378_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1163_c2_1dfb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_6ea6_return_output;
     -- n8_MUX[uxn_opcodes_h_l1182_c7_80b2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1182_c7_80b2_cond <= VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_cond;
     n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue;
     n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output := n8_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1182_c7_80b2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1182_c7_80b2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1182_c7_80b2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;

     -- MUX[uxn_opcodes_h_l1187_c21_9865] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1187_c21_9865_cond <= VAR_MUX_uxn_opcodes_h_l1187_c21_9865_cond;
     MUX_uxn_opcodes_h_l1187_c21_9865_iftrue <= VAR_MUX_uxn_opcodes_h_l1187_c21_9865_iftrue;
     MUX_uxn_opcodes_h_l1187_c21_9865_iffalse <= VAR_MUX_uxn_opcodes_h_l1187_c21_9865_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1187_c21_9865_return_output := MUX_uxn_opcodes_h_l1187_c21_9865_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1182_c7_80b2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;

     -- t8_MUX[uxn_opcodes_h_l1179_c7_4023] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1179_c7_4023_cond <= VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_cond;
     t8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue;
     t8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output := t8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue := VAR_MUX_uxn_opcodes_h_l1187_c21_9865_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1179_c7_4023] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;

     -- t8_MUX[uxn_opcodes_h_l1176_c7_04de] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1176_c7_04de_cond <= VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_cond;
     t8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue;
     t8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output := t8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1179_c7_4023] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1179_c7_4023] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1179_c7_4023] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;

     -- n8_MUX[uxn_opcodes_h_l1179_c7_4023] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1179_c7_4023_cond <= VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_cond;
     n8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue;
     n8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output := n8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1182_c7_80b2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_80b2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1176_c7_04de] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1176_c7_04de] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1176_c7_04de] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1179_c7_4023] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_return_output := result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;

     -- t8_MUX[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond <= VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond;
     t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue;
     t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output := t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1176_c7_04de] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;

     -- n8_MUX[uxn_opcodes_h_l1176_c7_04de] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1176_c7_04de_cond <= VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_cond;
     n8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue;
     n8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output := n8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_4023_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1176_c7_04de] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_return_output := result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;

     -- n8_MUX[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond <= VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond;
     n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue;
     n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output := n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_04de_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1163_c2_1dfb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output := result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1191_l1159_DUPLICATE_19d0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1191_l1159_DUPLICATE_19d0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_04b4(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_1dfb_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1191_l1159_DUPLICATE_19d0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l1191_l1159_DUPLICATE_19d0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
