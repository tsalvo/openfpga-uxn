-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity lth_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_6d7675a8;
architecture arch of lth_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2009_c6_1fc4]
signal BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2009_c1_1e91]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2009_c2_eac3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2009_c2_eac3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2009_c2_eac3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2009_c2_eac3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2009_c2_eac3]
signal result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2009_c2_eac3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2009_c2_eac3]
signal t8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2009_c2_eac3]
signal n8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2010_c3_ffb6[uxn_opcodes_h_l2010_c3_ffb6]
signal printf_uxn_opcodes_h_l2010_c3_ffb6_uxn_opcodes_h_l2010_c3_ffb6_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2014_c11_39d1]
signal BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2014_c7_152f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2014_c7_152f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2014_c7_152f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2014_c7_152f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2014_c7_152f]
signal result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2014_c7_152f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2014_c7_152f]
signal t8_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2014_c7_152f]
signal n8_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2017_c11_50bd]
signal BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2017_c7_2cb8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2017_c7_2cb8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2017_c7_2cb8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2017_c7_2cb8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2017_c7_2cb8]
signal result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2017_c7_2cb8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2017_c7_2cb8]
signal t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2017_c7_2cb8]
signal n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2021_c11_3eaa]
signal BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2021_c7_fa85]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2021_c7_fa85]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2021_c7_fa85]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2021_c7_fa85]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2021_c7_fa85]
signal result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2021_c7_fa85]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2021_c7_fa85]
signal n8_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2024_c11_29ca]
signal BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2024_c7_e18f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2024_c7_e18f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2024_c7_e18f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2024_c7_e18f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2024_c7_e18f]
signal result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2024_c7_e18f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2024_c7_e18f]
signal n8_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2027_c30_8c3c]
signal sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l2030_c21_f696]
signal BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2030_c21_206c]
signal MUX_uxn_opcodes_h_l2030_c21_206c_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2030_c21_206c_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2030_c21_206c_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2030_c21_206c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2032_c11_9e2a]
signal BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2032_c7_dcc9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2032_c7_dcc9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2032_c7_dcc9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4
BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_left,
BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_right,
BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3
result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3
result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3
result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3
result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output);

-- t8_MUX_uxn_opcodes_h_l2009_c2_eac3
t8_MUX_uxn_opcodes_h_l2009_c2_eac3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond,
t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue,
t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse,
t8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output);

-- n8_MUX_uxn_opcodes_h_l2009_c2_eac3
n8_MUX_uxn_opcodes_h_l2009_c2_eac3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond,
n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue,
n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse,
n8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output);

-- printf_uxn_opcodes_h_l2010_c3_ffb6_uxn_opcodes_h_l2010_c3_ffb6
printf_uxn_opcodes_h_l2010_c3_ffb6_uxn_opcodes_h_l2010_c3_ffb6 : entity work.printf_uxn_opcodes_h_l2010_c3_ffb6_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2010_c3_ffb6_uxn_opcodes_h_l2010_c3_ffb6_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1
BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_left,
BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_right,
BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f
result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f
result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f
result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f
result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output);

-- t8_MUX_uxn_opcodes_h_l2014_c7_152f
t8_MUX_uxn_opcodes_h_l2014_c7_152f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2014_c7_152f_cond,
t8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue,
t8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse,
t8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output);

-- n8_MUX_uxn_opcodes_h_l2014_c7_152f
n8_MUX_uxn_opcodes_h_l2014_c7_152f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2014_c7_152f_cond,
n8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue,
n8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse,
n8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd
BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_left,
BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_right,
BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8
result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8
result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8
result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8
result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output);

-- t8_MUX_uxn_opcodes_h_l2017_c7_2cb8
t8_MUX_uxn_opcodes_h_l2017_c7_2cb8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond,
t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue,
t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse,
t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output);

-- n8_MUX_uxn_opcodes_h_l2017_c7_2cb8
n8_MUX_uxn_opcodes_h_l2017_c7_2cb8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond,
n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue,
n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse,
n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa
BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_left,
BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_right,
BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85
result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85
result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85
result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85
result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_cond,
result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85
result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output);

-- n8_MUX_uxn_opcodes_h_l2021_c7_fa85
n8_MUX_uxn_opcodes_h_l2021_c7_fa85 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2021_c7_fa85_cond,
n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue,
n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse,
n8_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca
BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_left,
BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_right,
BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f
result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f
result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f
result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f
result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output);

-- n8_MUX_uxn_opcodes_h_l2024_c7_e18f
n8_MUX_uxn_opcodes_h_l2024_c7_e18f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2024_c7_e18f_cond,
n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue,
n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse,
n8_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c
sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_ins,
sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_x,
sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_y,
sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696
BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696 : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_left,
BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_right,
BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_return_output);

-- MUX_uxn_opcodes_h_l2030_c21_206c
MUX_uxn_opcodes_h_l2030_c21_206c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2030_c21_206c_cond,
MUX_uxn_opcodes_h_l2030_c21_206c_iftrue,
MUX_uxn_opcodes_h_l2030_c21_206c_iffalse,
MUX_uxn_opcodes_h_l2030_c21_206c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a
BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_left,
BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_right,
BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9
result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9
result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9
result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
 t8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
 n8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output,
 t8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output,
 n8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output,
 t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output,
 n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output,
 n8_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output,
 n8_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output,
 sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_return_output,
 BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_return_output,
 MUX_uxn_opcodes_h_l2030_c21_206c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2011_c3_f1b6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2010_c3_ffb6_uxn_opcodes_h_l2010_c3_ffb6_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2015_c3_1aa8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2019_c3_90cc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2022_c3_dccf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2029_c3_0914 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2024_c7_e18f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2030_c21_206c_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2030_c21_206c_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2030_c21_206c_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2030_c21_206c_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_b008_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_abcb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_64d0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_1efa_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2017_l2014_l2032_l2024_l2021_DUPLICATE_28bd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2038_l2005_DUPLICATE_c74b_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_opcodes_h_l2030_c21_206c_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2015_c3_1aa8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2015_c3_1aa8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2011_c3_f1b6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2011_c3_f1b6;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2029_c3_0914 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2029_c3_0914;
     VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2022_c3_dccf := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2022_c3_dccf;
     VAR_MUX_uxn_opcodes_h_l2030_c21_206c_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2019_c3_90cc := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2019_c3_90cc;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2014_c11_39d1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_b008 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_b008_return_output := result.is_sp_shift;

     -- BIN_OP_LT[uxn_opcodes_h_l2030_c21_f696] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_left;
     BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_return_output := BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2027_c30_8c3c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_ins;
     sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_x;
     sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_return_output := sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2024_c7_e18f] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2024_c7_e18f_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2032_c11_9e2a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2017_c11_50bd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2017_l2014_l2032_l2024_l2021_DUPLICATE_28bd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2017_l2014_l2032_l2024_l2021_DUPLICATE_28bd_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2021_c11_3eaa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_left;
     BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output := BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_abcb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_abcb_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2024_c11_29ca] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_left;
     BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output := BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_64d0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_64d0_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2009_c6_1fc4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_1efa LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_1efa_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2009_c6_1fc4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2014_c11_39d1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2017_c11_50bd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2021_c11_3eaa_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2024_c11_29ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2032_c11_9e2a_return_output;
     VAR_MUX_uxn_opcodes_h_l2030_c21_206c_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l2030_c21_f696_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_1efa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_1efa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_1efa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_1efa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_1efa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2017_l2014_l2032_l2024_l2021_DUPLICATE_28bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2017_l2014_l2032_l2024_l2021_DUPLICATE_28bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2017_l2014_l2032_l2024_l2021_DUPLICATE_28bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2017_l2014_l2032_l2024_l2021_DUPLICATE_28bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2017_l2014_l2032_l2024_l2021_DUPLICATE_28bd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_b008_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_b008_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_b008_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_b008_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_b008_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_abcb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_abcb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_abcb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_abcb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2032_l2021_DUPLICATE_abcb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_64d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_64d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_64d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_64d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2017_l2014_l2009_l2024_l2021_DUPLICATE_64d0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2024_c7_e18f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2027_c30_8c3c_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2032_c7_dcc9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output;

     -- n8_MUX[uxn_opcodes_h_l2024_c7_e18f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2024_c7_e18f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_cond;
     n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue;
     n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output := n8_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2009_c1_1e91] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2032_c7_dcc9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output;

     -- MUX[uxn_opcodes_h_l2030_c21_206c] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2030_c21_206c_cond <= VAR_MUX_uxn_opcodes_h_l2030_c21_206c_cond;
     MUX_uxn_opcodes_h_l2030_c21_206c_iftrue <= VAR_MUX_uxn_opcodes_h_l2030_c21_206c_iftrue;
     MUX_uxn_opcodes_h_l2030_c21_206c_iffalse <= VAR_MUX_uxn_opcodes_h_l2030_c21_206c_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2030_c21_206c_return_output := MUX_uxn_opcodes_h_l2030_c21_206c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2032_c7_dcc9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2024_c7_e18f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;

     -- t8_MUX[uxn_opcodes_h_l2017_c7_2cb8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond;
     t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue;
     t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output := t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2024_c7_e18f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue := VAR_MUX_uxn_opcodes_h_l2030_c21_206c_return_output;
     VAR_printf_uxn_opcodes_h_l2010_c3_ffb6_uxn_opcodes_h_l2010_c3_ffb6_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2009_c1_1e91_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2032_c7_dcc9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;
     -- n8_MUX[uxn_opcodes_h_l2021_c7_fa85] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2021_c7_fa85_cond <= VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_cond;
     n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue;
     n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output := n8_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2024_c7_e18f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2024_c7_e18f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2024_c7_e18f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;

     -- t8_MUX[uxn_opcodes_h_l2014_c7_152f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2014_c7_152f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_cond;
     t8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue;
     t8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output := t8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2021_c7_fa85] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2021_c7_fa85] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2024_c7_e18f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;

     -- printf_uxn_opcodes_h_l2010_c3_ffb6[uxn_opcodes_h_l2010_c3_ffb6] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2010_c3_ffb6_uxn_opcodes_h_l2010_c3_ffb6_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2010_c3_ffb6_uxn_opcodes_h_l2010_c3_ffb6_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2024_c7_e18f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2021_c7_fa85] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2017_c7_2cb8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2017_c7_2cb8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2021_c7_fa85] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output := result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;

     -- n8_MUX[uxn_opcodes_h_l2017_c7_2cb8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond;
     n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue;
     n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output := n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;

     -- t8_MUX[uxn_opcodes_h_l2009_c2_eac3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond <= VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond;
     t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue;
     t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output := t8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2021_c7_fa85] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2021_c7_fa85] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2021_c7_fa85_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2014_c7_152f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2017_c7_2cb8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2014_c7_152f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;

     -- n8_MUX[uxn_opcodes_h_l2014_c7_152f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2014_c7_152f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_cond;
     n8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue;
     n8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output := n8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2017_c7_2cb8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2017_c7_2cb8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2017_c7_2cb8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2017_c7_2cb8_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2009_c2_eac3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output;

     -- n8_MUX[uxn_opcodes_h_l2009_c2_eac3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond <= VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_cond;
     n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue;
     n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output := n8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2014_c7_152f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2014_c7_152f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2014_c7_152f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2014_c7_152f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2009_c2_eac3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2014_c7_152f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2009_c2_eac3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2009_c2_eac3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2009_c2_eac3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2009_c2_eac3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2038_l2005_DUPLICATE_c74b LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2038_l2005_DUPLICATE_c74b_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2009_c2_eac3_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2038_l2005_DUPLICATE_c74b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2038_l2005_DUPLICATE_c74b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
