-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity add_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end add_0CLK_f62d646e;
architecture arch of add_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l859_c6_6b3a]
signal BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l859_c1_f54f]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l859_c2_29f6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l859_c2_29f6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l859_c2_29f6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l859_c2_29f6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l859_c2_29f6]
signal result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l859_c2_29f6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l859_c2_29f6]
signal t8_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l859_c2_29f6]
signal n8_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l860_c3_41af[uxn_opcodes_h_l860_c3_41af]
signal printf_uxn_opcodes_h_l860_c3_41af_uxn_opcodes_h_l860_c3_41af_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l864_c11_df65]
signal BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l864_c7_261c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l864_c7_261c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l864_c7_261c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l864_c7_261c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l864_c7_261c]
signal result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l864_c7_261c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l864_c7_261c]
signal t8_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l864_c7_261c]
signal n8_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l867_c11_b6cc]
signal BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l867_c7_54d2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l867_c7_54d2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l867_c7_54d2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l867_c7_54d2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l867_c7_54d2]
signal result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l867_c7_54d2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l867_c7_54d2]
signal t8_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l867_c7_54d2]
signal n8_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l871_c11_50fe]
signal BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l871_c7_f41c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l871_c7_f41c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l871_c7_f41c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l871_c7_f41c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l871_c7_f41c]
signal result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l871_c7_f41c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l871_c7_f41c]
signal n8_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l874_c11_1e78]
signal BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l874_c7_32d7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l874_c7_32d7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l874_c7_32d7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l874_c7_32d7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l874_c7_32d7]
signal result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l874_c7_32d7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l874_c7_32d7]
signal n8_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l877_c30_20f8]
signal sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l880_c21_09cb]
signal BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_right : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l882_c11_ba38]
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l882_c7_2758]
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l882_c7_2758]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l882_c7_2758]
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a
BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_left,
BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_right,
BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6
result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6
result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6
result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_cond,
result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output);

-- t8_MUX_uxn_opcodes_h_l859_c2_29f6
t8_MUX_uxn_opcodes_h_l859_c2_29f6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l859_c2_29f6_cond,
t8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue,
t8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse,
t8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output);

-- n8_MUX_uxn_opcodes_h_l859_c2_29f6
n8_MUX_uxn_opcodes_h_l859_c2_29f6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l859_c2_29f6_cond,
n8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue,
n8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse,
n8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output);

-- printf_uxn_opcodes_h_l860_c3_41af_uxn_opcodes_h_l860_c3_41af
printf_uxn_opcodes_h_l860_c3_41af_uxn_opcodes_h_l860_c3_41af : entity work.printf_uxn_opcodes_h_l860_c3_41af_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l860_c3_41af_uxn_opcodes_h_l860_c3_41af_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65
BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_left,
BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_right,
BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c
result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c
result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c
result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c
result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_cond,
result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c
result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output);

-- t8_MUX_uxn_opcodes_h_l864_c7_261c
t8_MUX_uxn_opcodes_h_l864_c7_261c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l864_c7_261c_cond,
t8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue,
t8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse,
t8_MUX_uxn_opcodes_h_l864_c7_261c_return_output);

-- n8_MUX_uxn_opcodes_h_l864_c7_261c
n8_MUX_uxn_opcodes_h_l864_c7_261c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l864_c7_261c_cond,
n8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue,
n8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse,
n8_MUX_uxn_opcodes_h_l864_c7_261c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc
BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_left,
BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_right,
BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2
result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2
result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2
result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2
result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_cond,
result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2
result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output);

-- t8_MUX_uxn_opcodes_h_l867_c7_54d2
t8_MUX_uxn_opcodes_h_l867_c7_54d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l867_c7_54d2_cond,
t8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue,
t8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse,
t8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output);

-- n8_MUX_uxn_opcodes_h_l867_c7_54d2
n8_MUX_uxn_opcodes_h_l867_c7_54d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l867_c7_54d2_cond,
n8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue,
n8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse,
n8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe
BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_left,
BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_right,
BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c
result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c
result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c
result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c
result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_cond,
result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c
result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output);

-- n8_MUX_uxn_opcodes_h_l871_c7_f41c
n8_MUX_uxn_opcodes_h_l871_c7_f41c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l871_c7_f41c_cond,
n8_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue,
n8_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse,
n8_MUX_uxn_opcodes_h_l871_c7_f41c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78
BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_left,
BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_right,
BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7
result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7
result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7
result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7
result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_cond,
result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7
result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output);

-- n8_MUX_uxn_opcodes_h_l874_c7_32d7
n8_MUX_uxn_opcodes_h_l874_c7_32d7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l874_c7_32d7_cond,
n8_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue,
n8_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse,
n8_MUX_uxn_opcodes_h_l874_c7_32d7_return_output);

-- sp_relative_shift_uxn_opcodes_h_l877_c30_20f8
sp_relative_shift_uxn_opcodes_h_l877_c30_20f8 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_ins,
sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_x,
sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_y,
sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb
BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb : entity work.BIN_OP_PLUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_left,
BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_right,
BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38
BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_left,
BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_right,
BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
 t8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
 n8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output,
 t8_MUX_uxn_opcodes_h_l864_c7_261c_return_output,
 n8_MUX_uxn_opcodes_h_l864_c7_261c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output,
 t8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output,
 n8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output,
 n8_MUX_uxn_opcodes_h_l871_c7_f41c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output,
 n8_MUX_uxn_opcodes_h_l874_c7_32d7_return_output,
 sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l861_c3_6af8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l860_c3_41af_uxn_opcodes_h_l860_c3_41af_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l865_c3_11a8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l869_c3_37d1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l872_c3_a16b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_013a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l874_c7_32d7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l880_c3_c1a1 : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_a542_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_ff68_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_8b89_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_b872_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l864_l882_l874_l871_l867_DUPLICATE_0685_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l855_l888_DUPLICATE_42d0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l865_c3_11a8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l865_c3_11a8;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_013a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_013a;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l872_c3_a16b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l872_c3_a16b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l861_c3_6af8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l861_c3_6af8;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l869_c3_37d1 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l869_c3_37d1;
     VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iffalse := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l877_c30_20f8] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_ins;
     sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_x <= VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_x;
     sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_y <= VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_return_output := sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l874_c11_1e78] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_left;
     BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output := BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l874_c7_32d7] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l874_c7_32d7_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_ff68 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_ff68_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l864_c11_df65] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_left;
     BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output := BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_b872 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_b872_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l864_l882_l874_l871_l867_DUPLICATE_0685 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l864_l882_l874_l871_l867_DUPLICATE_0685_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l859_c6_6b3a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_left;
     BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output := BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l880_c21_09cb] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_left;
     BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_return_output := BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l867_c11_b6cc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_left;
     BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output := BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l882_c11_ba38] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_left;
     BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_return_output := BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_8b89 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_8b89_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l871_c11_50fe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_left;
     BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output := BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_a542 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_a542_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c6_6b3a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l864_c11_df65_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l867_c11_b6cc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l871_c11_50fe_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l874_c11_1e78_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_ba38_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l880_c3_c1a1 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l880_c21_09cb_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_b872_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_b872_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_b872_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_b872_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_b872_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l864_l882_l874_l871_l867_DUPLICATE_0685_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l864_l882_l874_l871_l867_DUPLICATE_0685_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l864_l882_l874_l871_l867_DUPLICATE_0685_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l864_l882_l874_l871_l867_DUPLICATE_0685_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l864_l882_l874_l871_l867_DUPLICATE_0685_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_a542_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_a542_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_a542_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_a542_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_a542_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_ff68_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_ff68_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_ff68_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_ff68_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l864_l859_l882_l871_l867_DUPLICATE_ff68_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_8b89_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_8b89_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_8b89_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_8b89_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l864_l859_l874_l871_l867_DUPLICATE_8b89_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l874_c7_32d7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l877_c30_20f8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue := VAR_result_u8_value_uxn_opcodes_h_l880_c3_c1a1;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l882_c7_2758] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l874_c7_32d7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l874_c7_32d7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_return_output := result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l882_c7_2758] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_return_output;

     -- n8_MUX[uxn_opcodes_h_l874_c7_32d7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l874_c7_32d7_cond <= VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_cond;
     n8_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue;
     n8_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_return_output := n8_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l882_c7_2758] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l859_c1_f54f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l874_c7_32d7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;

     -- t8_MUX[uxn_opcodes_h_l867_c7_54d2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l867_c7_54d2_cond <= VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_cond;
     t8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue;
     t8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output := t8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l860_c3_41af_uxn_opcodes_h_l860_c3_41af_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l859_c1_f54f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_2758_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_2758_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_2758_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;
     -- n8_MUX[uxn_opcodes_h_l871_c7_f41c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l871_c7_f41c_cond <= VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_cond;
     n8_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue;
     n8_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_return_output := n8_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l874_c7_32d7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;

     -- printf_uxn_opcodes_h_l860_c3_41af[uxn_opcodes_h_l860_c3_41af] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l860_c3_41af_uxn_opcodes_h_l860_c3_41af_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l860_c3_41af_uxn_opcodes_h_l860_c3_41af_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l871_c7_f41c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_return_output := result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;

     -- t8_MUX[uxn_opcodes_h_l864_c7_261c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l864_c7_261c_cond <= VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_cond;
     t8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue;
     t8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_return_output := t8_MUX_uxn_opcodes_h_l864_c7_261c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l871_c7_f41c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l874_c7_32d7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l874_c7_32d7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l871_c7_f41c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l874_c7_32d7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l864_c7_261c_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l867_c7_54d2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_return_output := result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l871_c7_f41c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l871_c7_f41c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l867_c7_54d2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;

     -- t8_MUX[uxn_opcodes_h_l859_c2_29f6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l859_c2_29f6_cond <= VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_cond;
     t8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue;
     t8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output := t8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output;

     -- n8_MUX[uxn_opcodes_h_l867_c7_54d2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l867_c7_54d2_cond <= VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_cond;
     n8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue;
     n8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output := n8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l871_c7_f41c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l867_c7_54d2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l871_c7_f41c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l867_c7_54d2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l864_c7_261c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_return_output := result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l867_c7_54d2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l864_c7_261c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l864_c7_261c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l867_c7_54d2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;

     -- n8_MUX[uxn_opcodes_h_l864_c7_261c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l864_c7_261c_cond <= VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_cond;
     n8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_iftrue;
     n8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_return_output := n8_MUX_uxn_opcodes_h_l864_c7_261c_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l864_c7_261c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l867_c7_54d2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l864_c7_261c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l864_c7_261c_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l859_c2_29f6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l864_c7_261c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l859_c2_29f6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_return_output := result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l864_c7_261c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l859_c2_29f6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output;

     -- n8_MUX[uxn_opcodes_h_l859_c2_29f6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l859_c2_29f6_cond <= VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_cond;
     n8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue;
     n8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output := n8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l864_c7_261c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l859_c2_29f6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l864_c7_261c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l864_c7_261c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l864_c7_261c_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l859_c2_29f6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l859_c2_29f6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l859_c2_29f6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l855_l888_DUPLICATE_42d0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l855_l888_DUPLICATE_42d0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c2_29f6_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c2_29f6_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l855_l888_DUPLICATE_42d0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l855_l888_DUPLICATE_42d0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
