-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity and_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end and_0CLK_f62d646e;
architecture arch of and_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l947_c6_4003]
signal BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l947_c1_0547]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l947_c2_05d6]
signal n8_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l947_c2_05d6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l947_c2_05d6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l947_c2_05d6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l947_c2_05d6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l947_c2_05d6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l947_c2_05d6]
signal result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l947_c2_05d6]
signal t8_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l948_c3_c3da[uxn_opcodes_h_l948_c3_c3da]
signal printf_uxn_opcodes_h_l948_c3_c3da_uxn_opcodes_h_l948_c3_c3da_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l952_c11_fac8]
signal BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l952_c7_8494]
signal n8_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l952_c7_8494]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l952_c7_8494]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l952_c7_8494]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l952_c7_8494]
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l952_c7_8494]
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l952_c7_8494]
signal result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l952_c7_8494]
signal t8_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l955_c11_6447]
signal BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l955_c7_39e5]
signal n8_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l955_c7_39e5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l955_c7_39e5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l955_c7_39e5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l955_c7_39e5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l955_c7_39e5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l955_c7_39e5]
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l955_c7_39e5]
signal t8_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l959_c11_db33]
signal BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l959_c7_fb24]
signal n8_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l959_c7_fb24]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l959_c7_fb24]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l959_c7_fb24]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l959_c7_fb24]
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l959_c7_fb24]
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l959_c7_fb24]
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l962_c11_e545]
signal BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l962_c7_d3ea]
signal n8_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l962_c7_d3ea]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l962_c7_d3ea]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l962_c7_d3ea]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l962_c7_d3ea]
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l962_c7_d3ea]
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l962_c7_d3ea]
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l965_c30_7635]
signal sp_relative_shift_uxn_opcodes_h_l965_c30_7635_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l965_c30_7635_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l965_c30_7635_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l965_c30_7635_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l968_c21_cb24]
signal BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l970_c11_ac9a]
signal BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l970_c7_7d3a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l970_c7_7d3a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l970_c7_7d3a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8cda( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003
BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_left,
BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_right,
BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_return_output);

-- n8_MUX_uxn_opcodes_h_l947_c2_05d6
n8_MUX_uxn_opcodes_h_l947_c2_05d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l947_c2_05d6_cond,
n8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue,
n8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse,
n8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6
result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6
result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6
result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6
result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6
result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_cond,
result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_return_output);

-- t8_MUX_uxn_opcodes_h_l947_c2_05d6
t8_MUX_uxn_opcodes_h_l947_c2_05d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l947_c2_05d6_cond,
t8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue,
t8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse,
t8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output);

-- printf_uxn_opcodes_h_l948_c3_c3da_uxn_opcodes_h_l948_c3_c3da
printf_uxn_opcodes_h_l948_c3_c3da_uxn_opcodes_h_l948_c3_c3da : entity work.printf_uxn_opcodes_h_l948_c3_c3da_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l948_c3_c3da_uxn_opcodes_h_l948_c3_c3da_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8
BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_left,
BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_right,
BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output);

-- n8_MUX_uxn_opcodes_h_l952_c7_8494
n8_MUX_uxn_opcodes_h_l952_c7_8494 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l952_c7_8494_cond,
n8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue,
n8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse,
n8_MUX_uxn_opcodes_h_l952_c7_8494_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494
result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494
result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494
result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_cond,
result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_return_output);

-- t8_MUX_uxn_opcodes_h_l952_c7_8494
t8_MUX_uxn_opcodes_h_l952_c7_8494 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l952_c7_8494_cond,
t8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue,
t8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse,
t8_MUX_uxn_opcodes_h_l952_c7_8494_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447
BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_left,
BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_right,
BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output);

-- n8_MUX_uxn_opcodes_h_l955_c7_39e5
n8_MUX_uxn_opcodes_h_l955_c7_39e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l955_c7_39e5_cond,
n8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue,
n8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse,
n8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5
result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_cond,
result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_return_output);

-- t8_MUX_uxn_opcodes_h_l955_c7_39e5
t8_MUX_uxn_opcodes_h_l955_c7_39e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l955_c7_39e5_cond,
t8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue,
t8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse,
t8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33
BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_left,
BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_right,
BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output);

-- n8_MUX_uxn_opcodes_h_l959_c7_fb24
n8_MUX_uxn_opcodes_h_l959_c7_fb24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l959_c7_fb24_cond,
n8_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue,
n8_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse,
n8_MUX_uxn_opcodes_h_l959_c7_fb24_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24
result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_cond,
result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545
BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_left,
BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_right,
BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output);

-- n8_MUX_uxn_opcodes_h_l962_c7_d3ea
n8_MUX_uxn_opcodes_h_l962_c7_d3ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l962_c7_d3ea_cond,
n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue,
n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse,
n8_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea
result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_cond,
result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output);

-- sp_relative_shift_uxn_opcodes_h_l965_c30_7635
sp_relative_shift_uxn_opcodes_h_l965_c30_7635 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l965_c30_7635_ins,
sp_relative_shift_uxn_opcodes_h_l965_c30_7635_x,
sp_relative_shift_uxn_opcodes_h_l965_c30_7635_y,
sp_relative_shift_uxn_opcodes_h_l965_c30_7635_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24
BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_left,
BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_right,
BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a
BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_left,
BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_right,
BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a
result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a
result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a
result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_return_output,
 n8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
 t8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output,
 n8_MUX_uxn_opcodes_h_l952_c7_8494_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_return_output,
 t8_MUX_uxn_opcodes_h_l952_c7_8494_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output,
 n8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_return_output,
 t8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output,
 n8_MUX_uxn_opcodes_h_l959_c7_fb24_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output,
 n8_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output,
 sp_relative_shift_uxn_opcodes_h_l965_c30_7635_return_output,
 BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l949_c3_b3cc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l948_c3_c3da_uxn_opcodes_h_l948_c3_c3da_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l953_c3_6662 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l957_c3_5ba9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l960_c3_b50f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l967_c3_5f8e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l962_c7_d3ea_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_229a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_b276_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_35f0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_e636_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l955_l952_l970_l962_l959_DUPLICATE_d8bf_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l976_l943_DUPLICATE_2e6c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l953_c3_6662 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l953_c3_6662;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l960_c3_b50f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l960_c3_b50f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l949_c3_b3cc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l949_c3_b3cc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l957_c3_5ba9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l957_c3_5ba9;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l967_c3_5f8e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l967_c3_5f8e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_right := to_unsigned(5, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_e636 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_e636_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_229a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_229a_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_35f0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_35f0_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l965_c30_7635] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l965_c30_7635_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_ins;
     sp_relative_shift_uxn_opcodes_h_l965_c30_7635_x <= VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_x;
     sp_relative_shift_uxn_opcodes_h_l965_c30_7635_y <= VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_return_output := sp_relative_shift_uxn_opcodes_h_l965_c30_7635_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l959_c11_db33] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_left;
     BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output := BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_b276 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_b276_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l955_l952_l970_l962_l959_DUPLICATE_d8bf LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l955_l952_l970_l962_l959_DUPLICATE_d8bf_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l955_c11_6447] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_left;
     BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output := BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l962_c11_e545] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_left;
     BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output := BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l970_c11_ac9a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_left;
     BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_return_output := BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l968_c21_cb24] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_left;
     BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_return_output := BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l952_c11_fac8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_left;
     BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output := BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l947_c6_4003] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_left;
     BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output := BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l962_c7_d3ea] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l962_c7_d3ea_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l968_c21_cb24_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l947_c6_4003_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l952_c11_fac8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_6447_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l959_c11_db33_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_e545_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l970_c11_ac9a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_229a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_229a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_229a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_229a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_229a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l955_l952_l970_l962_l959_DUPLICATE_d8bf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l955_l952_l970_l962_l959_DUPLICATE_d8bf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l955_l952_l970_l962_l959_DUPLICATE_d8bf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l955_l952_l970_l962_l959_DUPLICATE_d8bf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l955_l952_l970_l962_l959_DUPLICATE_d8bf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_b276_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_b276_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_b276_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_b276_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_b276_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_35f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_35f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_35f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_35f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l955_l952_l947_l970_l959_DUPLICATE_35f0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_e636_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_e636_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_e636_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_e636_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l955_l952_l947_l962_l959_DUPLICATE_e636_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l962_c7_d3ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l965_c30_7635_return_output;
     -- n8_MUX[uxn_opcodes_h_l962_c7_d3ea] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l962_c7_d3ea_cond <= VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_cond;
     n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue;
     n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output := n8_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l962_c7_d3ea] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l970_c7_7d3a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l947_c1_0547] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l962_c7_d3ea] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;

     -- t8_MUX[uxn_opcodes_h_l955_c7_39e5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l955_c7_39e5_cond <= VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_cond;
     t8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue;
     t8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output := t8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l970_c7_7d3a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l962_c7_d3ea] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_cond;
     result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output := result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l970_c7_7d3a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l948_c3_c3da_uxn_opcodes_h_l948_c3_c3da_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l947_c1_0547_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse := VAR_n8_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l970_c7_7d3a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse := VAR_t8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l959_c7_fb24] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_cond;
     result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_return_output := result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l962_c7_d3ea] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l962_c7_d3ea] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;

     -- printf_uxn_opcodes_h_l948_c3_c3da[uxn_opcodes_h_l948_c3_c3da] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l948_c3_c3da_uxn_opcodes_h_l948_c3_c3da_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l948_c3_c3da_uxn_opcodes_h_l948_c3_c3da_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_opc_done_MUX[uxn_opcodes_h_l962_c7_d3ea] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;

     -- t8_MUX[uxn_opcodes_h_l952_c7_8494] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l952_c7_8494_cond <= VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_cond;
     t8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue;
     t8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_return_output := t8_MUX_uxn_opcodes_h_l952_c7_8494_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l959_c7_fb24] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l959_c7_fb24] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;

     -- n8_MUX[uxn_opcodes_h_l959_c7_fb24] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l959_c7_fb24_cond <= VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_cond;
     n8_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue;
     n8_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_return_output := n8_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_d3ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l952_c7_8494_return_output;
     -- t8_MUX[uxn_opcodes_h_l947_c2_05d6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l947_c2_05d6_cond <= VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_cond;
     t8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue;
     t8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output := t8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output;

     -- n8_MUX[uxn_opcodes_h_l955_c7_39e5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l955_c7_39e5_cond <= VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_cond;
     n8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue;
     n8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output := n8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l959_c7_fb24] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l955_c7_39e5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l955_c7_39e5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l959_c7_fb24] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l955_c7_39e5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_return_output := result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l959_c7_fb24] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse := VAR_n8_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l959_c7_fb24_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l955_c7_39e5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l955_c7_39e5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l952_c7_8494] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_return_output;

     -- n8_MUX[uxn_opcodes_h_l952_c7_8494] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l952_c7_8494_cond <= VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_cond;
     n8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_iftrue;
     n8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_return_output := n8_MUX_uxn_opcodes_h_l952_c7_8494_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l955_c7_39e5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l952_c7_8494] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l952_c7_8494] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_cond;
     result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_return_output := result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l952_c7_8494_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_39e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l952_c7_8494_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l952_c7_8494_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l947_c2_05d6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_return_output := result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_return_output;

     -- n8_MUX[uxn_opcodes_h_l947_c2_05d6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l947_c2_05d6_cond <= VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_cond;
     n8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue;
     n8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output := n8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l952_c7_8494] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l947_c2_05d6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l952_c7_8494] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l952_c7_8494] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l947_c2_05d6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l947_c2_05d6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l952_c7_8494_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l952_c7_8494_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l952_c7_8494_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l947_c2_05d6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l947_c2_05d6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l947_c2_05d6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l976_l943_DUPLICATE_2e6c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l976_l943_DUPLICATE_2e6c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8cda(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l947_c2_05d6_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l947_c2_05d6_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l976_l943_DUPLICATE_2e6c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l976_l943_DUPLICATE_2e6c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
