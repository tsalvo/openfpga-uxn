-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 8
entity opc_dei2_0CLK_aa33bb56 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_dei2_0CLK_aa33bb56;
architecture arch of opc_dei2_0CLK_aa33bb56 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- t_register[uxn_opcodes_h_l707_c7_8d45]
signal t_register_uxn_opcodes_h_l707_c7_8d45_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_h_l707_c7_8d45_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_h_l707_c7_8d45_return_output : unsigned(7 downto 0);

-- set[uxn_opcodes_h_l708_c9_4ea8]
signal set_uxn_opcodes_h_l708_c9_4ea8_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_h_l708_c9_4ea8_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_h_l708_c9_4ea8_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_h_l708_c9_4ea8_k : unsigned(7 downto 0);
signal set_uxn_opcodes_h_l708_c9_4ea8_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_h_l708_c9_4ea8_add : signed(7 downto 0);
signal set_uxn_opcodes_h_l708_c9_4ea8_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l709_c6_51c3]
signal BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l710_c1_0a35]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_h_l709_c2_76f3]
signal result_MUX_uxn_opcodes_h_l709_c2_76f3_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_h_l709_c2_76f3_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_h_l709_c2_76f3_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_h_l709_c2_76f3_return_output : unsigned(0 downto 0);

-- dei[uxn_opcodes_h_l711_c3_06eb]
signal dei_uxn_opcodes_h_l711_c3_06eb_CLOCK_ENABLE : unsigned(0 downto 0);
signal dei_uxn_opcodes_h_l711_c3_06eb_stack_index : unsigned(0 downto 0);
signal dei_uxn_opcodes_h_l711_c3_06eb_stack_offset : unsigned(7 downto 0);
signal dei_uxn_opcodes_h_l711_c3_06eb_addr : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l712_c23_41bd]
signal BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_return_output : unsigned(8 downto 0);

-- dei[uxn_opcodes_h_l712_c3_c77b]
signal dei_uxn_opcodes_h_l712_c3_c77b_CLOCK_ENABLE : unsigned(0 downto 0);
signal dei_uxn_opcodes_h_l712_c3_c77b_stack_index : unsigned(0 downto 0);
signal dei_uxn_opcodes_h_l712_c3_c77b_stack_offset : unsigned(7 downto 0);
signal dei_uxn_opcodes_h_l712_c3_c77b_addr : unsigned(7 downto 0);


begin

-- SUBMODULE INSTANCES 
-- t_register_uxn_opcodes_h_l707_c7_8d45
t_register_uxn_opcodes_h_l707_c7_8d45 : entity work.t_register_0CLK_0e5af5c0 port map (
clk,
t_register_uxn_opcodes_h_l707_c7_8d45_CLOCK_ENABLE,
t_register_uxn_opcodes_h_l707_c7_8d45_stack_index,
t_register_uxn_opcodes_h_l707_c7_8d45_return_output);

-- set_uxn_opcodes_h_l708_c9_4ea8
set_uxn_opcodes_h_l708_c9_4ea8 : entity work.set_0CLK_082cb698 port map (
clk,
set_uxn_opcodes_h_l708_c9_4ea8_CLOCK_ENABLE,
set_uxn_opcodes_h_l708_c9_4ea8_stack_index,
set_uxn_opcodes_h_l708_c9_4ea8_ins,
set_uxn_opcodes_h_l708_c9_4ea8_k,
set_uxn_opcodes_h_l708_c9_4ea8_mul,
set_uxn_opcodes_h_l708_c9_4ea8_add,
set_uxn_opcodes_h_l708_c9_4ea8_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3
BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_left,
BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_right,
BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_return_output);

-- result_MUX_uxn_opcodes_h_l709_c2_76f3
result_MUX_uxn_opcodes_h_l709_c2_76f3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_h_l709_c2_76f3_cond,
result_MUX_uxn_opcodes_h_l709_c2_76f3_iftrue,
result_MUX_uxn_opcodes_h_l709_c2_76f3_iffalse,
result_MUX_uxn_opcodes_h_l709_c2_76f3_return_output);

-- dei_uxn_opcodes_h_l711_c3_06eb
dei_uxn_opcodes_h_l711_c3_06eb : entity work.dei_0CLK_f8b40cb1 port map (
clk,
dei_uxn_opcodes_h_l711_c3_06eb_CLOCK_ENABLE,
dei_uxn_opcodes_h_l711_c3_06eb_stack_index,
dei_uxn_opcodes_h_l711_c3_06eb_stack_offset,
dei_uxn_opcodes_h_l711_c3_06eb_addr);

-- BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd
BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_left,
BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_right,
BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_return_output);

-- dei_uxn_opcodes_h_l712_c3_c77b
dei_uxn_opcodes_h_l712_c3_c77b : entity work.dei_0CLK_f8b40cb1 port map (
clk,
dei_uxn_opcodes_h_l712_c3_c77b_CLOCK_ENABLE,
dei_uxn_opcodes_h_l712_c3_c77b_stack_index,
dei_uxn_opcodes_h_l712_c3_c77b_stack_offset,
dei_uxn_opcodes_h_l712_c3_c77b_addr);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 stack_index,
 ins,
 k,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 t_register_uxn_opcodes_h_l707_c7_8d45_return_output,
 set_uxn_opcodes_h_l708_c9_4ea8_return_output,
 BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_return_output,
 result_MUX_uxn_opcodes_h_l709_c2_76f3_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_h_l707_c7_8d45_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_h_l707_c7_8d45_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_h_l707_c7_8d45_return_output : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_h_l708_c9_4ea8_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_h_l708_c9_4ea8_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_h_l708_c9_4ea8_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_h_l708_c9_4ea8_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_h_l708_c9_4ea8_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_h_l708_c9_4ea8_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_h_l708_c9_4ea8_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_cond : unsigned(0 downto 0);
 variable VAR_dei_uxn_opcodes_h_l711_c3_06eb_stack_index : unsigned(0 downto 0);
 variable VAR_dei_uxn_opcodes_h_l711_c3_06eb_stack_offset : unsigned(7 downto 0);
 variable VAR_dei_uxn_opcodes_h_l711_c3_06eb_addr : unsigned(7 downto 0);
 variable VAR_dei_uxn_opcodes_h_l711_c3_06eb_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_dei_uxn_opcodes_h_l712_c3_c77b_stack_index : unsigned(0 downto 0);
 variable VAR_dei_uxn_opcodes_h_l712_c3_c77b_stack_offset : unsigned(7 downto 0);
 variable VAR_dei_uxn_opcodes_h_l712_c3_c77b_addr : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_return_output : unsigned(8 downto 0);
 variable VAR_dei_uxn_opcodes_h_l712_c3_c77b_CLOCK_ENABLE : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_iffalse := to_unsigned(0, 1);
     VAR_dei_uxn_opcodes_h_l712_c3_c77b_stack_offset := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_right := to_unsigned(1, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iftrue := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_h_l708_c9_4ea8_mul := resize(to_unsigned(1, 1), 8);
     VAR_set_uxn_opcodes_h_l708_c9_4ea8_add := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_right := to_unsigned(0, 1);
     VAR_dei_uxn_opcodes_h_l711_c3_06eb_stack_offset := resize(to_unsigned(1, 1), 8);
     VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iffalse := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_h_l708_c9_4ea8_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_t_register_uxn_opcodes_h_l707_c7_8d45_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_h_l708_c9_4ea8_ins := VAR_ins;
     VAR_set_uxn_opcodes_h_l708_c9_4ea8_k := VAR_k;
     VAR_dei_uxn_opcodes_h_l711_c3_06eb_stack_index := VAR_stack_index;
     VAR_dei_uxn_opcodes_h_l712_c3_c77b_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_h_l708_c9_4ea8_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_h_l707_c7_8d45_stack_index := VAR_stack_index;
     -- t_register[uxn_opcodes_h_l707_c7_8d45] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_h_l707_c7_8d45_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_h_l707_c7_8d45_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_h_l707_c7_8d45_stack_index <= VAR_t_register_uxn_opcodes_h_l707_c7_8d45_stack_index;
     -- Outputs
     VAR_t_register_uxn_opcodes_h_l707_c7_8d45_return_output := t_register_uxn_opcodes_h_l707_c7_8d45_return_output;

     -- set[uxn_opcodes_h_l708_c9_4ea8] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_h_l708_c9_4ea8_CLOCK_ENABLE <= VAR_set_uxn_opcodes_h_l708_c9_4ea8_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_h_l708_c9_4ea8_stack_index <= VAR_set_uxn_opcodes_h_l708_c9_4ea8_stack_index;
     set_uxn_opcodes_h_l708_c9_4ea8_ins <= VAR_set_uxn_opcodes_h_l708_c9_4ea8_ins;
     set_uxn_opcodes_h_l708_c9_4ea8_k <= VAR_set_uxn_opcodes_h_l708_c9_4ea8_k;
     set_uxn_opcodes_h_l708_c9_4ea8_mul <= VAR_set_uxn_opcodes_h_l708_c9_4ea8_mul;
     set_uxn_opcodes_h_l708_c9_4ea8_add <= VAR_set_uxn_opcodes_h_l708_c9_4ea8_add;
     -- Outputs
     VAR_set_uxn_opcodes_h_l708_c9_4ea8_return_output := set_uxn_opcodes_h_l708_c9_4ea8_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_left := VAR_set_uxn_opcodes_h_l708_c9_4ea8_return_output;
     REG_VAR_tmp8 := VAR_set_uxn_opcodes_h_l708_c9_4ea8_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_left := VAR_t_register_uxn_opcodes_h_l707_c7_8d45_return_output;
     VAR_dei_uxn_opcodes_h_l711_c3_06eb_addr := VAR_t_register_uxn_opcodes_h_l707_c7_8d45_return_output;
     REG_VAR_t8 := VAR_t_register_uxn_opcodes_h_l707_c7_8d45_return_output;
     -- BIN_OP_PLUS[uxn_opcodes_h_l712_c23_41bd] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_left;
     BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_return_output := BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l709_c6_51c3] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_left;
     BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_return_output := BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_return_output;
     VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l709_c6_51c3_return_output;
     VAR_dei_uxn_opcodes_h_l712_c3_c77b_addr := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l712_c23_41bd_return_output, 8);
     -- result_MUX[uxn_opcodes_h_l709_c2_76f3] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_h_l709_c2_76f3_cond <= VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_cond;
     result_MUX_uxn_opcodes_h_l709_c2_76f3_iftrue <= VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_iftrue;
     result_MUX_uxn_opcodes_h_l709_c2_76f3_iffalse <= VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_return_output := result_MUX_uxn_opcodes_h_l709_c2_76f3_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l710_c1_0a35] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_return_output;

     -- Submodule level 3
     VAR_dei_uxn_opcodes_h_l711_c3_06eb_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_return_output;
     VAR_dei_uxn_opcodes_h_l712_c3_c77b_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l710_c1_0a35_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_h_l709_c2_76f3_return_output;
     -- dei[uxn_opcodes_h_l712_c3_c77b] LATENCY=0
     -- Clock enable
     dei_uxn_opcodes_h_l712_c3_c77b_CLOCK_ENABLE <= VAR_dei_uxn_opcodes_h_l712_c3_c77b_CLOCK_ENABLE;
     -- Inputs
     dei_uxn_opcodes_h_l712_c3_c77b_stack_index <= VAR_dei_uxn_opcodes_h_l712_c3_c77b_stack_index;
     dei_uxn_opcodes_h_l712_c3_c77b_stack_offset <= VAR_dei_uxn_opcodes_h_l712_c3_c77b_stack_offset;
     dei_uxn_opcodes_h_l712_c3_c77b_addr <= VAR_dei_uxn_opcodes_h_l712_c3_c77b_addr;
     -- Outputs

     -- dei[uxn_opcodes_h_l711_c3_06eb] LATENCY=0
     -- Clock enable
     dei_uxn_opcodes_h_l711_c3_06eb_CLOCK_ENABLE <= VAR_dei_uxn_opcodes_h_l711_c3_06eb_CLOCK_ENABLE;
     -- Inputs
     dei_uxn_opcodes_h_l711_c3_06eb_stack_index <= VAR_dei_uxn_opcodes_h_l711_c3_06eb_stack_index;
     dei_uxn_opcodes_h_l711_c3_06eb_stack_offset <= VAR_dei_uxn_opcodes_h_l711_c3_06eb_stack_offset;
     dei_uxn_opcodes_h_l711_c3_06eb_addr <= VAR_dei_uxn_opcodes_h_l711_c3_06eb_addr;
     -- Outputs

     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
