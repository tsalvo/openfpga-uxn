-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 33
entity VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28 is
port(
 elem_val : in unsigned(7 downto 0);
 ref_toks_0 : in uint8_t_16;
 var_dim_0 : in unsigned(3 downto 0);
 return_output : out uint8_t_array_16_t);
end VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28;
architecture arch of VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iftrue : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iffalse : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iftrue : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iffalse : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iftrue : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iffalse : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_return_output : unsigned(0 downto 0);

-- rv_data_13_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03]
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_cond : unsigned(0 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iftrue : unsigned(7 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iffalse : unsigned(7 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_return_output : unsigned(0 downto 0);

-- rv_data_10_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75]
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_cond : unsigned(0 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iftrue : unsigned(7 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iffalse : unsigned(7 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iftrue : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iffalse : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iftrue : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iffalse : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_return_output : unsigned(0 downto 0);

-- rv_data_11_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef]
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_cond : unsigned(0 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iftrue : unsigned(7 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iffalse : unsigned(7 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_return_output : unsigned(0 downto 0);

-- rv_data_8_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17]
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_cond : unsigned(0 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iftrue : unsigned(7 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iffalse : unsigned(7 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_return_output : unsigned(0 downto 0);

-- rv_data_14_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8]
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_cond : unsigned(0 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iftrue : unsigned(7 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iffalse : unsigned(7 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iftrue : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iffalse : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iftrue : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iffalse : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iftrue : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iffalse : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_return_output : unsigned(0 downto 0);

-- rv_data_9_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251]
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_cond : unsigned(0 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iftrue : unsigned(7 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iffalse : unsigned(7 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_return_output : unsigned(0 downto 0);

-- rv_data_12_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007]
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_cond : unsigned(0 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iftrue : unsigned(7 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iffalse : unsigned(7 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_return_output : unsigned(0 downto 0);

-- rv_data_15_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42]
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_cond : unsigned(0 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iftrue : unsigned(7 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iffalse : unsigned(7 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_return_output : unsigned(7 downto 0);

function CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_8c3c( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint8_t_array_16_t is
 
  variable base : uint8_t_array_16_t; 
  variable return_output : uint8_t_array_16_t;
begin
      base.data(4) := ref_toks_0;
      base.data(1) := ref_toks_1;
      base.data(7) := ref_toks_2;
      base.data(13) := ref_toks_3;
      base.data(10) := ref_toks_4;
      base.data(2) := ref_toks_5;
      base.data(5) := ref_toks_6;
      base.data(11) := ref_toks_7;
      base.data(8) := ref_toks_8;
      base.data(14) := ref_toks_9;
      base.data(0) := ref_toks_10;
      base.data(6) := ref_toks_11;
      base.data(3) := ref_toks_12;
      base.data(9) := ref_toks_13;
      base.data(12) := ref_toks_14;
      base.data(15) := ref_toks_15;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_return_output);

-- rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_cond,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iftrue,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iffalse,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_return_output);

-- rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_cond,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iftrue,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iffalse,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_return_output);

-- rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_cond,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iftrue,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iffalse,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_return_output);

-- rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_cond,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iftrue,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iffalse,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_return_output);

-- rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_cond,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iftrue,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iffalse,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_return_output);

-- rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_cond,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iftrue,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iffalse,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_return_output);

-- rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_cond,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iftrue,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iffalse,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_return_output);

-- rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_cond,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iftrue,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iffalse,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_return_output,
 rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_return_output,
 rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_return_output,
 rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_return_output,
 rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_return_output,
 rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_return_output,
 rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_return_output,
 rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_return_output,
 rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(7 downto 0);
 variable VAR_ref_toks_0 : uint8_t_16;
 variable VAR_var_dim_0 : unsigned(3 downto 0);
 variable VAR_return_output : uint8_t_array_16_t;
 variable VAR_base : uint8_t_16;
 variable VAR_rv : uint8_t_array_16_t;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_4b72_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_4685_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_6728_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_fb4a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_6ffb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_a17f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_c37e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c16_271a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_4d33_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_f317_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c15_640a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_eb42_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_e579_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_4099_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_dc47_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_b8f8_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_8c3c_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_0f58_return_output : uint8_t_array_16_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_right := to_unsigned(15, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_right := to_unsigned(9, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_right := to_unsigned(13, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_right := to_unsigned(10, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_right := to_unsigned(11, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_right := to_unsigned(8, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_right := to_unsigned(14, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_right := to_unsigned(12, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_right := to_unsigned(5, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iftrue := VAR_elem_val;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iftrue := VAR_elem_val;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iftrue := VAR_elem_val;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iftrue := VAR_elem_val;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iftrue := VAR_elem_val;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iftrue := VAR_elem_val;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iftrue := VAR_elem_val;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iftrue := VAR_elem_val;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_left := VAR_var_dim_0;
     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_4_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_4b72] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_4b72_return_output := VAR_ref_toks_0(4);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_7_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_6728] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_6728_return_output := VAR_ref_toks_0(7);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_13_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_fb4a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_fb4a_return_output := VAR_ref_toks_0(13);

     -- CONST_REF_RD_uint8_t_uint8_t_16_8_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_4d33] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_4d33_return_output := VAR_ref_toks_0(8);

     -- CONST_REF_RD_uint8_t_uint8_t_16_14_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_f317] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_f317_return_output := VAR_ref_toks_0(14);

     -- CONST_REF_RD_uint8_t_uint8_t_16_1_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_4685] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_4685_return_output := VAR_ref_toks_0(1);

     -- CONST_REF_RD_uint8_t_uint8_t_16_11_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c16_271a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c16_271a_return_output := VAR_ref_toks_0(11);

     -- CONST_REF_RD_uint8_t_uint8_t_16_15_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_b8f8] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_b8f8_return_output := VAR_ref_toks_0(15);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_9_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_4099] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_4099_return_output := VAR_ref_toks_0(9);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_0_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c15_640a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c15_640a_return_output := VAR_ref_toks_0(0);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_6_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_eb42] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_eb42_return_output := VAR_ref_toks_0(6);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_5_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_c37e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_c37e_return_output := VAR_ref_toks_0(5);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_10_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_6ffb] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_6ffb_return_output := VAR_ref_toks_0(10);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_2_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_a17f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_a17f_return_output := VAR_ref_toks_0(2);

     -- CONST_REF_RD_uint8_t_uint8_t_16_3_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_e579] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_e579_return_output := VAR_ref_toks_0(3);

     -- CONST_REF_RD_uint8_t_uint8_t_16_12_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_dc47] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_dc47_return_output := VAR_ref_toks_0(12);

     -- Submodule level 1
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_e3c5_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_992d_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_1fd1_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_e2a1_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_8fff_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_9058_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_ced8_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_fb81_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_29f0_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_c846_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_b73f_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_470c_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_d52d_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ab_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_f63b_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_f702_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c15_640a_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_6ffb_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c16_271a_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c16_dc47_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_fb4a_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_f317_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_b8f8_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_4685_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_a17f_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_e579_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_4b72_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_c37e_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_eb42_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_6728_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_4d33_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_4099_return_output;
     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84] LATENCY=0
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_iffalse;
     -- Outputs
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_return_output;

     -- rv_data_14_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8] LATENCY=0
     -- Inputs
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_cond <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_cond;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iftrue <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iftrue;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iffalse <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_iffalse;
     -- Outputs
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_return_output := rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_return_output;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9] LATENCY=0
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_iffalse;
     -- Outputs
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_return_output;

     -- rv_data_15_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42] LATENCY=0
     -- Inputs
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_cond <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_cond;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iftrue <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iftrue;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iffalse <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_iffalse;
     -- Outputs
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_return_output := rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_return_output;

     -- rv_data_9_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251] LATENCY=0
     -- Inputs
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_cond <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_cond;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iftrue <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iftrue;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iffalse <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_iffalse;
     -- Outputs
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_return_output := rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_return_output;

     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398] LATENCY=0
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_iffalse;
     -- Outputs
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_return_output;

     -- rv_data_8_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17] LATENCY=0
     -- Inputs
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_cond <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_cond;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iftrue <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iftrue;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iffalse <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_iffalse;
     -- Outputs
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_return_output := rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_return_output;

     -- rv_data_13_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03] LATENCY=0
     -- Inputs
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_cond <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_cond;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iftrue <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iftrue;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iffalse <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_iffalse;
     -- Outputs
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_return_output := rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_return_output;

     -- rv_data_10_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75] LATENCY=0
     -- Inputs
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_cond <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_cond;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iftrue <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iftrue;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iffalse <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_iffalse;
     -- Outputs
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_return_output := rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_return_output;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4] LATENCY=0
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_iffalse;
     -- Outputs
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_return_output;

     -- rv_data_11_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef] LATENCY=0
     -- Inputs
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_cond <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_cond;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iftrue <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iftrue;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iffalse <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_iffalse;
     -- Outputs
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_return_output := rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_return_output;

     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d] LATENCY=0
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_iffalse;
     -- Outputs
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_return_output;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548] LATENCY=0
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_iffalse;
     -- Outputs
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_return_output;

     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98] LATENCY=0
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_iffalse;
     -- Outputs
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_return_output;

     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6] LATENCY=0
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_iffalse;
     -- Outputs
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_return_output;

     -- rv_data_12_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007] LATENCY=0
     -- Inputs
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_cond <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_cond;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iftrue <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iftrue;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iffalse <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_iffalse;
     -- Outputs
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_return_output := rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_return_output;

     -- Submodule level 2
     -- CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_8c3c[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_0f58] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_8c3c_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_0f58_return_output := CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_8c3c(
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_a398_return_output,
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d84_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_96b4_return_output,
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_ea03_return_output,
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_ee75_return_output,
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_b8d6_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_c21d_return_output,
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_b6ef_return_output,
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_8b17_return_output,
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0cd8_return_output,
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_3548_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6a98_return_output,
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_aac9_return_output,
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_5251_return_output,
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_8007_return_output,
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_ec42_return_output);

     -- Submodule level 3
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_8c3c_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_0f58_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
