-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity dei_0CLK_99af4b2a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 controller0_buttons : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dei_0CLK_99af4b2a;
architecture arch of dei_0CLK_99af4b2a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal has_written_to_t : unsigned(0 downto 0) := to_unsigned(0, 1);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal device_in_result : device_in_result_t := device_in_result_t_NULL;
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_has_written_to_t : unsigned(0 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_device_in_result : device_in_result_t;
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l403_c6_c3fc]
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l419_c7_c017]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l403_c2_13cb]
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l403_c2_13cb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l403_c2_13cb]
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l403_c2_13cb]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l403_c2_13cb]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l403_c2_13cb]
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(7 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l403_c2_13cb]
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l403_c2_13cb]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l403_c2_13cb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l403_c2_13cb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l403_c2_13cb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(3 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l403_c2_13cb]
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l403_c2_13cb]
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : device_in_result_t;

-- t8_MUX[uxn_opcodes_h_l403_c2_13cb]
signal t8_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l419_c11_25cb]
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l422_c1_9a11]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l419_c7_c017]
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l419_c7_c017]
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l419_c7_c017]
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l419_c7_c017]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l419_c7_c017]
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l419_c7_c017]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(3 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l419_c7_c017]
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l419_c7_c017]
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_return_output : device_in_result_t;

-- t8_MUX[uxn_opcodes_h_l419_c7_c017]
signal t8_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l420_c30_166a]
signal sp_relative_shift_uxn_opcodes_h_l420_c30_166a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_166a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_166a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l420_c30_166a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l424_c9_0934]
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l424_c9_b813]
signal MUX_uxn_opcodes_h_l424_c9_b813_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_b813_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_b813_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l424_c9_b813_return_output : unsigned(7 downto 0);

-- UNARY_OP_NOT[uxn_opcodes_h_l425_c8_28c5]
signal UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l425_c1_f56d]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l425_c3_ce36]
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l425_c3_ce36]
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l425_c3_ce36]
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l425_c3_ce36]
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l425_c3_ce36]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(3 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l425_c3_ce36]
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l425_c3_ce36]
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : device_in_result_t;

-- BIN_OP_MINUS[uxn_opcodes_h_l426_c37_7448]
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_right : unsigned(1 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_return_output : unsigned(7 downto 0);

-- device_in[uxn_opcodes_h_l426_c23_f255]
signal device_in_uxn_opcodes_h_l426_c23_f255_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_f255_device_address : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_f255_phase : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_f255_controller0_buttons : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_f255_previous_device_ram_read : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l426_c23_f255_return_output : device_in_result_t;

-- UNARY_OP_NOT[uxn_opcodes_h_l429_c9_2390]
signal UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l429_c4_2961]
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l429_c4_2961]
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l429_c4_2961]
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l429_c4_2961]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_return_output : unsigned(3 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l429_c4_2961]
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_return_output : unsigned(0 downto 0);

function CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6( ref_toks_0 : device_in_result_t;
 ref_toks_1 : unsigned) return device_in_result_t is
 
  variable base : device_in_result_t; 
  variable return_output : device_in_result_t;
begin
      base := ref_toks_0;
      base.is_dei_done := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_76ef( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : signed;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_device_ram_write := ref_toks_4;
      base.is_pc_updated := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.device_ram_address := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.sp_relative_shift := ref_toks_9;
      base.is_opc_done := ref_toks_10;
      base.stack_address_sp_offset := ref_toks_11;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc
BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_left,
BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_right,
BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb
result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb
device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- t8_MUX_uxn_opcodes_h_l403_c2_13cb
t8_MUX_uxn_opcodes_h_l403_c2_13cb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l403_c2_13cb_cond,
t8_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue,
t8_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse,
t8_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb
BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_left,
BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_right,
BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017
result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_cond,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_cond,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l419_c7_c017
device_in_result_MUX_uxn_opcodes_h_l419_c7_c017 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_cond,
device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iftrue,
device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iffalse,
device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_return_output);

-- t8_MUX_uxn_opcodes_h_l419_c7_c017
t8_MUX_uxn_opcodes_h_l419_c7_c017 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l419_c7_c017_cond,
t8_MUX_uxn_opcodes_h_l419_c7_c017_iftrue,
t8_MUX_uxn_opcodes_h_l419_c7_c017_iffalse,
t8_MUX_uxn_opcodes_h_l419_c7_c017_return_output);

-- sp_relative_shift_uxn_opcodes_h_l420_c30_166a
sp_relative_shift_uxn_opcodes_h_l420_c30_166a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l420_c30_166a_ins,
sp_relative_shift_uxn_opcodes_h_l420_c30_166a_x,
sp_relative_shift_uxn_opcodes_h_l420_c30_166a_y,
sp_relative_shift_uxn_opcodes_h_l420_c30_166a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934
BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_left,
BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_right,
BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_return_output);

-- MUX_uxn_opcodes_h_l424_c9_b813
MUX_uxn_opcodes_h_l424_c9_b813 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l424_c9_b813_cond,
MUX_uxn_opcodes_h_l424_c9_b813_iftrue,
MUX_uxn_opcodes_h_l424_c9_b813_iffalse,
MUX_uxn_opcodes_h_l424_c9_b813_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_expr,
UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36
result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_cond,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_cond,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36
device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_cond,
device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue,
device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse,
device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448 : entity work.BIN_OP_MINUS_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_left,
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_right,
BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_return_output);

-- device_in_uxn_opcodes_h_l426_c23_f255
device_in_uxn_opcodes_h_l426_c23_f255 : entity work.device_in_0CLK_50065acf port map (
clk,
device_in_uxn_opcodes_h_l426_c23_f255_CLOCK_ENABLE,
device_in_uxn_opcodes_h_l426_c23_f255_device_address,
device_in_uxn_opcodes_h_l426_c23_f255_phase,
device_in_uxn_opcodes_h_l426_c23_f255_controller0_buttons,
device_in_uxn_opcodes_h_l426_c23_f255_previous_device_ram_read,
device_in_uxn_opcodes_h_l426_c23_f255_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_expr,
UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961
result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_cond,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_cond,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 controller0_buttons,
 previous_stack_read,
 previous_device_ram_read,
 -- Registers
 has_written_to_t,
 t8,
 device_in_result,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 t8_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_return_output,
 device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_return_output,
 t8_MUX_uxn_opcodes_h_l419_c7_c017_return_output,
 sp_relative_shift_uxn_opcodes_h_l420_c30_166a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_return_output,
 MUX_uxn_opcodes_h_l424_c9_b813_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_return_output,
 device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_return_output,
 device_in_uxn_opcodes_h_l426_c23_f255_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_controller0_buttons : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_e8da : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_8637 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : device_in_result_t;
 variable VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_13cb_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_41aa : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_b813_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_b813_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_b813_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l424_c9_b813_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_1d16_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iffalse : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_cond : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_f255_device_address : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_f255_phase : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_f255_controller0_buttons : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_f255_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_return_output : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_f255_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l426_c23_f255_return_output : device_in_result_t;
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_8cc4_return_output : unsigned(7 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_5154 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_cond : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_fc6c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l419_l403_l425_l429_DUPLICATE_2165_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l419_l403_l425_DUPLICATE_9cab_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_9897_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_d7b6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_a105_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_76ef_uxn_opcodes_h_l441_l397_DUPLICATE_d0ed_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_has_written_to_t : unsigned(0 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_device_in_result : device_in_result_t;
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_has_written_to_t := has_written_to_t;
  REG_VAR_t8 := t8;
  REG_VAR_device_in_result := device_in_result;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_right := to_unsigned(0, 1);
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iftrue := to_unsigned(0, 1);
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_8637 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l414_c3_8637;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_5154 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l431_c5_5154;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iffalse := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_right := to_unsigned(2, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_right := to_unsigned(2, 2);
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_e8da := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l408_c3_e8da;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_41aa := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iffalse := VAR_result_sp_relative_shift_uxn_opcodes_h_l423_c3_41aa;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_controller0_buttons := controller0_buttons;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iffalse := VAR_CLOCK_ENABLE;
     VAR_device_in_uxn_opcodes_h_l426_c23_f255_controller0_buttons := VAR_controller0_buttons;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iftrue := device_in_result;
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse := device_in_result;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_expr := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iffalse := has_written_to_t;
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_left := VAR_phase;
     VAR_device_in_uxn_opcodes_h_l426_c23_f255_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_MUX_uxn_opcodes_h_l424_c9_b813_iftrue := VAR_previous_stack_read;
     VAR_MUX_uxn_opcodes_h_l424_c9_b813_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_iftrue := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_9897 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_9897_return_output := result.is_opc_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_13cb_return_output := result.is_vram_write;

     -- UNARY_OP_NOT[uxn_opcodes_h_l429_c9_2390] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_return_output := UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l403_c6_c3fc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_left;
     BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output := BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;

     -- CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d[uxn_opcodes_h_l432_c23_fc6c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_fc6c_return_output := device_in_result.dei_value;

     -- sp_relative_shift[uxn_opcodes_h_l420_c30_166a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l420_c30_166a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_ins;
     sp_relative_shift_uxn_opcodes_h_l420_c30_166a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_x;
     sp_relative_shift_uxn_opcodes_h_l420_c30_166a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_return_output := sp_relative_shift_uxn_opcodes_h_l420_c30_166a_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_a105 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_a105_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l419_c11_25cb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_left;
     BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output := BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output;

     -- result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_13cb_return_output := result.is_device_ram_write;

     -- device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_13cb_return_output := CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6(
     device_in_result,
     to_unsigned(0, 1));

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l419_l403_l425_DUPLICATE_9cab LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l419_l403_l425_DUPLICATE_9cab_return_output := result.device_ram_address;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_13cb_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l419_l403_l425_l429_DUPLICATE_2165 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l419_l403_l425_l429_DUPLICATE_2165_return_output := result.u8_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_13cb_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d[uxn_opcodes_h_l425_c8_1d16] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_1d16_return_output := device_in_result.is_dei_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l424_c9_0934] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_left;
     BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_return_output := BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_13cb_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_d7b6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_d7b6_return_output := result.is_stack_write;

     -- BIN_OP_MINUS[uxn_opcodes_h_l426_c37_7448] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_left;
     BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_return_output := BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l403_c6_c3fc_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l419_c11_25cb_return_output;
     VAR_MUX_uxn_opcodes_h_l424_c9_b813_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c9_0934_return_output;
     VAR_device_in_uxn_opcodes_h_l426_c23_f255_phase := VAR_BIN_OP_MINUS_uxn_opcodes_h_l426_c37_7448_return_output;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_expr := VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l425_c8_1d16_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_9897_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_9897_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_9897_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_d7b6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l419_l425_DUPLICATE_d7b6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_a105_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_a105_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l419_l425_l429_DUPLICATE_a105_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l432_c23_fc6c_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l419_l403_l425_DUPLICATE_9cab_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l419_l403_l425_DUPLICATE_9cab_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l419_l403_l425_DUPLICATE_9cab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l419_l403_l425_l429_DUPLICATE_2165_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l419_l403_l425_l429_DUPLICATE_2165_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l419_l403_l425_l429_DUPLICATE_2165_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l419_l403_l425_l429_DUPLICATE_2165_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l429_c9_2390_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue := VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l403_c2_13cb_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l403_c2_13cb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l403_c2_13cb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l403_c2_13cb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l403_c2_13cb_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l403_c2_13cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l420_c30_166a_return_output;
     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l429_c4_2961] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_cond;
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_return_output := result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_return_output;

     -- UNARY_OP_NOT[uxn_opcodes_h_l425_c8_28c5] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output := UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l429_c4_2961] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_return_output := has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l429_c4_2961] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l419_c7_c017] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- MUX[uxn_opcodes_h_l424_c9_b813] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l424_c9_b813_cond <= VAR_MUX_uxn_opcodes_h_l424_c9_b813_cond;
     MUX_uxn_opcodes_h_l424_c9_b813_iftrue <= VAR_MUX_uxn_opcodes_h_l424_c9_b813_iftrue;
     MUX_uxn_opcodes_h_l424_c9_b813_iffalse <= VAR_MUX_uxn_opcodes_h_l424_c9_b813_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l424_c9_b813_return_output := MUX_uxn_opcodes_h_l424_c9_b813_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l429_c4_2961] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l429_c4_2961] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l419_c7_c017] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l419_c7_c017_return_output;
     VAR_device_in_uxn_opcodes_h_l426_c23_f255_device_address := VAR_MUX_uxn_opcodes_h_l424_c9_b813_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_iffalse := VAR_MUX_uxn_opcodes_h_l424_c9_b813_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l425_c8_28c5_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l429_c4_2961_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l429_c4_2961_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l429_c4_2961_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l419_c7_c017_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l429_c4_2961_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l429_c4_2961_return_output;
     -- t8_MUX[uxn_opcodes_h_l419_c7_c017] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l419_c7_c017_cond <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_cond;
     t8_MUX_uxn_opcodes_h_l419_c7_c017_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_iftrue;
     t8_MUX_uxn_opcodes_h_l419_c7_c017_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_return_output := t8_MUX_uxn_opcodes_h_l419_c7_c017_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l425_c3_ce36] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l425_c3_ce36] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_return_output := has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l425_c3_ce36] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l422_c1_9a11] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l425_c3_ce36] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_cond;
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_return_output := result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l425_c3_ce36] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;

     -- Submodule level 3
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l422_c1_9a11_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_t8_MUX_uxn_opcodes_h_l419_c7_c017_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l425_c1_f56d] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_return_output;

     -- t8_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     t8_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     t8_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := t8_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l419_c7_c017] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l419_c7_c017] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l419_c7_c017] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_return_output := has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l419_c7_c017] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_cond;
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_return_output := result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l419_c7_c017] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_return_output;

     -- Submodule level 4
     VAR_device_in_uxn_opcodes_h_l426_c23_f255_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l425_c1_f56d_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l419_c7_c017_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l419_c7_c017_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l419_c7_c017_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l419_c7_c017_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l419_c7_c017_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;
     -- device_in[uxn_opcodes_h_l426_c23_f255] LATENCY=0
     -- Clock enable
     device_in_uxn_opcodes_h_l426_c23_f255_CLOCK_ENABLE <= VAR_device_in_uxn_opcodes_h_l426_c23_f255_CLOCK_ENABLE;
     -- Inputs
     device_in_uxn_opcodes_h_l426_c23_f255_device_address <= VAR_device_in_uxn_opcodes_h_l426_c23_f255_device_address;
     device_in_uxn_opcodes_h_l426_c23_f255_phase <= VAR_device_in_uxn_opcodes_h_l426_c23_f255_phase;
     device_in_uxn_opcodes_h_l426_c23_f255_controller0_buttons <= VAR_device_in_uxn_opcodes_h_l426_c23_f255_controller0_buttons;
     device_in_uxn_opcodes_h_l426_c23_f255_previous_device_ram_read <= VAR_device_in_uxn_opcodes_h_l426_c23_f255_previous_device_ram_read;
     -- Outputs
     VAR_device_in_uxn_opcodes_h_l426_c23_f255_return_output := device_in_uxn_opcodes_h_l426_c23_f255_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- Submodule level 5
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue := VAR_device_in_uxn_opcodes_h_l426_c23_f255_return_output;
     REG_VAR_has_written_to_t := VAR_has_written_to_t_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;
     -- CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d[uxn_opcodes_h_l427_c32_8cc4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_8cc4_return_output := VAR_device_in_uxn_opcodes_h_l426_c23_f255_return_output.device_ram_address;

     -- device_in_result_MUX[uxn_opcodes_h_l425_c3_ce36] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_cond;
     device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_return_output := device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;

     -- Submodule level 6
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l427_c32_8cc4_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;
     -- device_in_result_MUX[uxn_opcodes_h_l419_c7_c017] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_cond;
     device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_return_output := device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l425_c3_ce36] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;

     -- Submodule level 7
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l419_c7_c017_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l425_c3_ce36_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l419_c7_c017] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_return_output;

     -- device_in_result_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- Submodule level 8
     REG_VAR_device_in_result := VAR_device_in_result_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l419_c7_c017_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l403_c2_13cb] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_76ef_uxn_opcodes_h_l441_l397_DUPLICATE_d0ed LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_76ef_uxn_opcodes_h_l441_l397_DUPLICATE_d0ed_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_76ef(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l403_c2_13cb_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l403_c2_13cb_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_76ef_uxn_opcodes_h_l441_l397_DUPLICATE_d0ed_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_76ef_uxn_opcodes_h_l441_l397_DUPLICATE_d0ed_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_has_written_to_t <= REG_VAR_has_written_to_t;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_device_in_result <= REG_VAR_device_in_result;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     has_written_to_t <= REG_COMB_has_written_to_t;
     t8 <= REG_COMB_t8;
     device_in_result <= REG_COMB_device_in_result;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
