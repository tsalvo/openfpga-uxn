-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity rot_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_b288bfb7;
architecture arch of rot_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2639_c6_b9bb]
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2639_c2_3b6f]
signal t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2652_c11_a7b9]
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2652_c7_3ed9]
signal l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2652_c7_3ed9]
signal n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2652_c7_3ed9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2652_c7_3ed9]
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2652_c7_3ed9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2652_c7_3ed9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2652_c7_3ed9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2652_c7_3ed9]
signal t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2655_c11_409d]
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2655_c7_8cfa]
signal l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2655_c7_8cfa]
signal n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2655_c7_8cfa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2655_c7_8cfa]
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2655_c7_8cfa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2655_c7_8cfa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2655_c7_8cfa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2655_c7_8cfa]
signal t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2659_c11_387a]
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2659_c7_037b]
signal l8_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2659_c7_037b]
signal n8_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2659_c7_037b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2659_c7_037b]
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2659_c7_037b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2659_c7_037b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2659_c7_037b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2661_c30_8a74]
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2666_c11_9521]
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2666_c7_8d7e]
signal l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2666_c7_8d7e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2666_c7_8d7e]
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2666_c7_8d7e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2666_c7_8d7e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_7531]
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_7ca7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_7ca7]
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_7ca7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_b856( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_left,
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_right,
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output);

-- l8_MUX_uxn_opcodes_h_l2639_c2_3b6f
l8_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- n8_MUX_uxn_opcodes_h_l2639_c2_3b6f
n8_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- t8_MUX_uxn_opcodes_h_l2639_c2_3b6f
t8_MUX_uxn_opcodes_h_l2639_c2_3b6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond,
t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue,
t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse,
t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_left,
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_right,
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output);

-- l8_MUX_uxn_opcodes_h_l2652_c7_3ed9
l8_MUX_uxn_opcodes_h_l2652_c7_3ed9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond,
l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue,
l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse,
l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output);

-- n8_MUX_uxn_opcodes_h_l2652_c7_3ed9
n8_MUX_uxn_opcodes_h_l2652_c7_3ed9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond,
n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue,
n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse,
n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output);

-- t8_MUX_uxn_opcodes_h_l2652_c7_3ed9
t8_MUX_uxn_opcodes_h_l2652_c7_3ed9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond,
t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue,
t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse,
t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_left,
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_right,
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output);

-- l8_MUX_uxn_opcodes_h_l2655_c7_8cfa
l8_MUX_uxn_opcodes_h_l2655_c7_8cfa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond,
l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue,
l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse,
l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output);

-- n8_MUX_uxn_opcodes_h_l2655_c7_8cfa
n8_MUX_uxn_opcodes_h_l2655_c7_8cfa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond,
n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue,
n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse,
n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output);

-- t8_MUX_uxn_opcodes_h_l2655_c7_8cfa
t8_MUX_uxn_opcodes_h_l2655_c7_8cfa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond,
t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue,
t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse,
t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_left,
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_right,
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output);

-- l8_MUX_uxn_opcodes_h_l2659_c7_037b
l8_MUX_uxn_opcodes_h_l2659_c7_037b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2659_c7_037b_cond,
l8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue,
l8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse,
l8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output);

-- n8_MUX_uxn_opcodes_h_l2659_c7_037b
n8_MUX_uxn_opcodes_h_l2659_c7_037b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2659_c7_037b_cond,
n8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue,
n8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse,
n8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74
sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_ins,
sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_x,
sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_y,
sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_left,
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_right,
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_return_output);

-- l8_MUX_uxn_opcodes_h_l2666_c7_8d7e
l8_MUX_uxn_opcodes_h_l2666_c7_8d7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond,
l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue,
l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse,
l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_left,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_right,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output,
 l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output,
 l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output,
 n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output,
 t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output,
 l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output,
 n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output,
 t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output,
 l8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output,
 n8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_return_output,
 sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_return_output,
 l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_0d0b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_c488 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_b165 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_1d62 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_6fff : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_a940 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_b5ec : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_435e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_7ca7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2639_l2672_l2652_DUPLICATE_fe35_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_cfc3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2666_l2652_DUPLICATE_3fed_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_e925_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2678_l2635_DUPLICATE_4dfa_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_b165 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_b165;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_right := to_unsigned(5, 3);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_c488 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_c488;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_1d62 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_1d62;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_a940 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_a940;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_435e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_435e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_right := to_unsigned(4, 3);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_b5ec := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_b5ec;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_0d0b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_0d0b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_6fff := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_6fff;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2666_l2652_DUPLICATE_3fed LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2666_l2652_DUPLICATE_3fed_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2659_c11_387a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_e925 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_e925_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2639_l2672_l2652_DUPLICATE_fe35 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2639_l2672_l2652_DUPLICATE_fe35_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2652_c11_a7b9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output := result.is_pc_updated;

     -- sp_relative_shift[uxn_opcodes_h_l2661_c30_8a74] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_ins;
     sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_x;
     sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_return_output := sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2666_c11_9521] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_left;
     BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_return_output := BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2672_c7_7ca7] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_7ca7_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2639_c6_b9bb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2655_c11_409d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_7531] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_left;
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_return_output := BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_cfc3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_cfc3_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_b9bb_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_a7b9_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_409d_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_387a_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_9521_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_7531_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2666_l2652_DUPLICATE_3fed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2666_l2652_DUPLICATE_3fed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2666_l2652_DUPLICATE_3fed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_e925_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_e925_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_e925_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_e925_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2659_l2655_l2652_l2672_l2666_DUPLICATE_e925_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_cfc3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_cfc3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_cfc3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2639_l2672_l2652_DUPLICATE_fe35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2639_l2672_l2652_DUPLICATE_fe35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2639_l2672_l2652_DUPLICATE_fe35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2639_l2672_l2652_DUPLICATE_fe35_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_3b6f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_7ca7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_8a74_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_7ca7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output;

     -- t8_MUX[uxn_opcodes_h_l2655_c7_8cfa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond;
     t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue;
     t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output := t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2666_c7_8d7e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output;

     -- l8_MUX[uxn_opcodes_h_l2666_c7_8d7e] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond;
     l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue;
     l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output := l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_7ca7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2659_c7_037b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;

     -- n8_MUX[uxn_opcodes_h_l2659_c7_037b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2659_c7_037b_cond <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_cond;
     n8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue;
     n8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output := n8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_7ca7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_7ca7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2655_c7_8cfa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2659_c7_037b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2666_c7_8d7e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2655_c7_8cfa] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond;
     n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue;
     n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output := n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2666_c7_8d7e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output;

     -- t8_MUX[uxn_opcodes_h_l2652_c7_3ed9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond;
     t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue;
     t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output := t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2666_c7_8d7e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output;

     -- l8_MUX[uxn_opcodes_h_l2659_c7_037b] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2659_c7_037b_cond <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_cond;
     l8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue;
     l8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output := l8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_8d7e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2659_c7_037b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2659_c7_037b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2655_c7_8cfa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;

     -- t8_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2659_c7_037b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;

     -- l8_MUX[uxn_opcodes_h_l2655_c7_8cfa] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond;
     l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue;
     l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output := l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;

     -- n8_MUX[uxn_opcodes_h_l2652_c7_3ed9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond;
     n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue;
     n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output := n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2652_c7_3ed9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_037b_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2655_c7_8cfa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2655_c7_8cfa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output := result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2652_c7_3ed9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2655_c7_8cfa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;

     -- n8_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- l8_MUX[uxn_opcodes_h_l2652_c7_3ed9] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond;
     l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue;
     l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output := l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_8cfa_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2652_c7_3ed9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;

     -- l8_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2652_c7_3ed9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2652_c7_3ed9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_3ed9_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c2_3b6f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2678_l2635_DUPLICATE_4dfa LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2678_l2635_DUPLICATE_4dfa_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_b856(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_3b6f_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2678_l2635_DUPLICATE_4dfa_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2678_l2635_DUPLICATE_4dfa_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
