-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity sub_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub_0CLK_64d180f1;
architecture arch of sub_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2484_c6_f294]
signal BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2484_c2_62f2]
signal t8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2484_c2_62f2]
signal n8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2484_c2_62f2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2484_c2_62f2]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2484_c2_62f2]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2484_c2_62f2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2484_c2_62f2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2484_c2_62f2]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2484_c2_62f2]
signal result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2484_c2_62f2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2484_c2_62f2]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2497_c11_5887]
signal BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2497_c7_a179]
signal t8_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2497_c7_a179]
signal n8_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2497_c7_a179]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2497_c7_a179]
signal result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2497_c7_a179]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2497_c7_a179]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2497_c7_a179]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2500_c11_bc9d]
signal BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2500_c7_c64a]
signal t8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2500_c7_c64a]
signal n8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2500_c7_c64a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2500_c7_c64a]
signal result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2500_c7_c64a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2500_c7_c64a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2500_c7_c64a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2503_c11_4f33]
signal BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2503_c7_01c0]
signal n8_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2503_c7_01c0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2503_c7_01c0]
signal result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2503_c7_01c0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2503_c7_01c0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2503_c7_01c0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2505_c30_9cc4]
signal sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2508_c21_8823]
signal BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294
BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_left,
BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_right,
BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output);

-- t8_MUX_uxn_opcodes_h_l2484_c2_62f2
t8_MUX_uxn_opcodes_h_l2484_c2_62f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond,
t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue,
t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse,
t8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

-- n8_MUX_uxn_opcodes_h_l2484_c2_62f2
n8_MUX_uxn_opcodes_h_l2484_c2_62f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond,
n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue,
n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse,
n8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2
result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2
result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2
result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2
result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2
result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2
result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887
BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_left,
BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_right,
BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output);

-- t8_MUX_uxn_opcodes_h_l2497_c7_a179
t8_MUX_uxn_opcodes_h_l2497_c7_a179 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2497_c7_a179_cond,
t8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue,
t8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse,
t8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output);

-- n8_MUX_uxn_opcodes_h_l2497_c7_a179
n8_MUX_uxn_opcodes_h_l2497_c7_a179 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2497_c7_a179_cond,
n8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue,
n8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse,
n8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179
result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179
result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_cond,
result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179
result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179
result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d
BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_left,
BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_right,
BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output);

-- t8_MUX_uxn_opcodes_h_l2500_c7_c64a
t8_MUX_uxn_opcodes_h_l2500_c7_c64a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond,
t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue,
t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse,
t8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output);

-- n8_MUX_uxn_opcodes_h_l2500_c7_c64a
n8_MUX_uxn_opcodes_h_l2500_c7_c64a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond,
n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue,
n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse,
n8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a
result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a
result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a
result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33
BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_left,
BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_right,
BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output);

-- n8_MUX_uxn_opcodes_h_l2503_c7_01c0
n8_MUX_uxn_opcodes_h_l2503_c7_01c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2503_c7_01c0_cond,
n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue,
n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse,
n8_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0
result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0
result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0
result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4
sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_ins,
sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_x,
sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_y,
sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823
BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_left,
BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_right,
BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output,
 t8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
 n8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output,
 t8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output,
 n8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output,
 t8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output,
 n8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output,
 n8_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output,
 sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2489_c3_e7ac : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2494_c3_d9ca : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2498_c3_a4bd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2507_c3_cbf9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2500_l2484_l2503_l2497_DUPLICATE_ab54_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_6dcc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_be1e_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_73a4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2500_l2503_DUPLICATE_5d0c_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2512_l2480_DUPLICATE_2d89_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_right := to_unsigned(3, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2489_c3_e7ac := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2489_c3_e7ac;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2507_c3_cbf9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2507_c3_cbf9;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2494_c3_d9ca := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2494_c3_d9ca;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2498_c3_a4bd := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2498_c3_a4bd;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_6dcc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_6dcc_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2500_l2503_DUPLICATE_5d0c LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2500_l2503_DUPLICATE_5d0c_return_output := result.stack_address_sp_offset;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2508_c21_8823] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2500_l2484_l2503_l2497_DUPLICATE_ab54 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2500_l2484_l2503_l2497_DUPLICATE_ab54_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2503_c11_4f33] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_left;
     BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output := BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2497_c11_5887] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_left;
     BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output := BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2484_c6_f294] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_left;
     BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output := BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2505_c30_9cc4] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_ins;
     sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_x;
     sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_return_output := sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_73a4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_73a4_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output := result.is_ram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_be1e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_be1e_return_output := result.sp_relative_shift;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2500_c11_bc9d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output := result.is_stack_index_flipped;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2484_c6_f294_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_5887_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2500_c11_bc9d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2503_c11_4f33_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2508_c21_8823_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_be1e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_be1e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_be1e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_6dcc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_6dcc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_6dcc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_73a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_73a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2500_l2503_l2497_DUPLICATE_73a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2500_l2503_DUPLICATE_5d0c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2500_l2503_DUPLICATE_5d0c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2500_l2484_l2503_l2497_DUPLICATE_ab54_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2500_l2484_l2503_l2497_DUPLICATE_ab54_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2500_l2484_l2503_l2497_DUPLICATE_ab54_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2500_l2484_l2503_l2497_DUPLICATE_ab54_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2484_c2_62f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2505_c30_9cc4_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2503_c7_01c0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2503_c7_01c0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;

     -- t8_MUX[uxn_opcodes_h_l2500_c7_c64a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond <= VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond;
     t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue;
     t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output := t8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;

     -- n8_MUX[uxn_opcodes_h_l2503_c7_01c0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2503_c7_01c0_cond <= VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_cond;
     n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue;
     n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output := n8_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2503_c7_01c0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2503_c7_01c0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2503_c7_01c0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2503_c7_01c0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2500_c7_c64a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2500_c7_c64a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;

     -- t8_MUX[uxn_opcodes_h_l2497_c7_a179] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2497_c7_a179_cond <= VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_cond;
     t8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue;
     t8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output := t8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2500_c7_c64a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2500_c7_c64a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2500_c7_c64a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;

     -- n8_MUX[uxn_opcodes_h_l2500_c7_c64a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_cond;
     n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iftrue;
     n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output := n8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2500_c7_c64a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2497_c7_a179] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2497_c7_a179] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;

     -- n8_MUX[uxn_opcodes_h_l2497_c7_a179] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2497_c7_a179_cond <= VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_cond;
     n8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue;
     n8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output := n8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;

     -- t8_MUX[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond <= VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond;
     t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue;
     t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output := t8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2497_c7_a179] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2497_c7_a179] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2497_c7_a179] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_return_output := result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_a179_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;
     -- n8_MUX[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond <= VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_cond;
     n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue;
     n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output := n8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2484_c2_62f2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2512_l2480_DUPLICATE_2d89 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2512_l2480_DUPLICATE_2d89_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2484_c2_62f2_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2512_l2480_DUPLICATE_2d89_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2512_l2480_DUPLICATE_2d89_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
