-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity neq_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_226c8821;
architecture arch of neq_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1259_c6_fc5d]
signal BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1259_c2_3184]
signal n8_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1259_c2_3184]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1259_c2_3184]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1259_c2_3184]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1259_c2_3184]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1259_c2_3184]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1259_c2_3184]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1259_c2_3184]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1259_c2_3184]
signal result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1259_c2_3184]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1259_c2_3184]
signal t8_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1272_c11_ef64]
signal BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1272_c7_0c0a]
signal n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1272_c7_0c0a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1272_c7_0c0a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1272_c7_0c0a]
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1272_c7_0c0a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1272_c7_0c0a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1272_c7_0c0a]
signal t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1275_c11_4299]
signal BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1275_c7_1e59]
signal n8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1275_c7_1e59]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1275_c7_1e59]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1275_c7_1e59]
signal result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1275_c7_1e59]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1275_c7_1e59]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1275_c7_1e59]
signal t8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1278_c11_d4fe]
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1278_c7_ea66]
signal n8_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1278_c7_ea66]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1278_c7_ea66]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1278_c7_ea66]
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1278_c7_ea66]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1278_c7_ea66]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1280_c30_37ba]
signal sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1283_c21_0bcf]
signal BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1283_c21_0ea6]
signal MUX_uxn_opcodes_h_l1283_c21_0ea6_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1283_c21_0ea6_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1283_c21_0ea6_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1283_c21_0ea6_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a47b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d
BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_left,
BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_right,
BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output);

-- n8_MUX_uxn_opcodes_h_l1259_c2_3184
n8_MUX_uxn_opcodes_h_l1259_c2_3184 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1259_c2_3184_cond,
n8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue,
n8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse,
n8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184
result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184
result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184
result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184
result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184
result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184
result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_cond,
result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184
result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

-- t8_MUX_uxn_opcodes_h_l1259_c2_3184
t8_MUX_uxn_opcodes_h_l1259_c2_3184 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1259_c2_3184_cond,
t8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue,
t8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse,
t8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_left,
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_right,
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output);

-- n8_MUX_uxn_opcodes_h_l1272_c7_0c0a
n8_MUX_uxn_opcodes_h_l1272_c7_0c0a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond,
n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue,
n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse,
n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output);

-- t8_MUX_uxn_opcodes_h_l1272_c7_0c0a
t8_MUX_uxn_opcodes_h_l1272_c7_0c0a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond,
t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue,
t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse,
t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299
BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_left,
BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_right,
BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output);

-- n8_MUX_uxn_opcodes_h_l1275_c7_1e59
n8_MUX_uxn_opcodes_h_l1275_c7_1e59 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond,
n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue,
n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse,
n8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59
result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59
result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59
result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_cond,
result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59
result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output);

-- t8_MUX_uxn_opcodes_h_l1275_c7_1e59
t8_MUX_uxn_opcodes_h_l1275_c7_1e59 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond,
t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue,
t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse,
t8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_left,
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_right,
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output);

-- n8_MUX_uxn_opcodes_h_l1278_c7_ea66
n8_MUX_uxn_opcodes_h_l1278_c7_ea66 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1278_c7_ea66_cond,
n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue,
n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse,
n8_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_cond,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba
sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_ins,
sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_x,
sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_y,
sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf
BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_left,
BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_right,
BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_return_output);

-- MUX_uxn_opcodes_h_l1283_c21_0ea6
MUX_uxn_opcodes_h_l1283_c21_0ea6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1283_c21_0ea6_cond,
MUX_uxn_opcodes_h_l1283_c21_0ea6_iftrue,
MUX_uxn_opcodes_h_l1283_c21_0ea6_iffalse,
MUX_uxn_opcodes_h_l1283_c21_0ea6_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output,
 n8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
 t8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output,
 n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output,
 t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output,
 n8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output,
 t8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output,
 n8_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output,
 sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_return_output,
 MUX_uxn_opcodes_h_l1283_c21_0ea6_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1264_c3_eca4 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1269_c3_d97e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1273_c3_0f76 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1282_c3_9ccd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_b3b5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_a811_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_5f50_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_947c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1275_l1278_DUPLICATE_e823_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1287_l1255_DUPLICATE_5dcc_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1273_c3_0f76 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1273_c3_0f76;
     VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1269_c3_d97e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1269_c3_d97e;
     VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1264_c3_eca4 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1264_c3_eca4;
     VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1282_c3_9ccd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1282_c3_9ccd;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_right := to_unsigned(3, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse := t8;
     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1259_c2_3184_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1272_c11_ef64] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_left;
     BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output := BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_5f50 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_5f50_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_947c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_947c_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1275_c11_4299] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_left;
     BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output := BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1259_c2_3184_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1275_l1278_DUPLICATE_e823 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1275_l1278_DUPLICATE_e823_return_output := result.stack_address_sp_offset;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1259_c2_3184_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1278_c11_d4fe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_left;
     BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output := BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_a811 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_a811_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_b3b5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_b3b5_return_output := result.u8_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1259_c2_3184_return_output := result.is_pc_updated;

     -- sp_relative_shift[uxn_opcodes_h_l1280_c30_37ba] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_ins;
     sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_x;
     sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_return_output := sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1259_c6_fc5d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1283_c21_0bcf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_left;
     BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_return_output := BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_fc5d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_ef64_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_4299_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_d4fe_return_output;
     VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_0bcf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_5f50_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_5f50_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_5f50_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_a811_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_a811_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_a811_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_947c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_947c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_947c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1275_l1278_DUPLICATE_e823_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1275_l1278_DUPLICATE_e823_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_b3b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_b3b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_b3b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_b3b5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1259_c2_3184_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1259_c2_3184_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1259_c2_3184_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1259_c2_3184_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_37ba_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1278_c7_ea66] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;

     -- t8_MUX[uxn_opcodes_h_l1275_c7_1e59] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond <= VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond;
     t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue;
     t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output := t8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1278_c7_ea66] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1278_c7_ea66] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;

     -- n8_MUX[uxn_opcodes_h_l1278_c7_ea66] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1278_c7_ea66_cond <= VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_cond;
     n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue;
     n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output := n8_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1278_c7_ea66] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;

     -- MUX[uxn_opcodes_h_l1283_c21_0ea6] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1283_c21_0ea6_cond <= VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_cond;
     MUX_uxn_opcodes_h_l1283_c21_0ea6_iftrue <= VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_iftrue;
     MUX_uxn_opcodes_h_l1283_c21_0ea6_iffalse <= VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_return_output := MUX_uxn_opcodes_h_l1283_c21_0ea6_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue := VAR_MUX_uxn_opcodes_h_l1283_c21_0ea6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1275_c7_1e59] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1275_c7_1e59] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;

     -- t8_MUX[uxn_opcodes_h_l1272_c7_0c0a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond;
     t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue;
     t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output := t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1278_c7_ea66] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output := result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;

     -- n8_MUX[uxn_opcodes_h_l1275_c7_1e59] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond <= VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_cond;
     n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue;
     n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output := n8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1275_c7_1e59] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1275_c7_1e59] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_ea66_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1275_c7_1e59] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output := result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1272_c7_0c0a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1272_c7_0c0a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;

     -- n8_MUX[uxn_opcodes_h_l1272_c7_0c0a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond;
     n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue;
     n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output := n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;

     -- t8_MUX[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1259_c2_3184_cond <= VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_cond;
     t8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue;
     t8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output := t8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1272_c7_0c0a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1272_c7_0c0a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_1e59_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;
     -- n8_MUX[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1259_c2_3184_cond <= VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_cond;
     n8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue;
     n8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output := n8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1272_c7_0c0a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_0c0a_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1259_c2_3184] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_return_output := result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1287_l1255_DUPLICATE_5dcc LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1287_l1255_DUPLICATE_5dcc_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a47b(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_3184_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_3184_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1287_l1255_DUPLICATE_5dcc_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1287_l1255_DUPLICATE_5dcc_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
