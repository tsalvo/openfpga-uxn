-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity sub_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub_0CLK_64d180f1;
architecture arch of sub_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2478_c6_46ee]
signal BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2478_c2_8fc1]
signal t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2478_c2_8fc1]
signal n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2478_c2_8fc1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2478_c2_8fc1]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2478_c2_8fc1]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2478_c2_8fc1]
signal result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2478_c2_8fc1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2478_c2_8fc1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2478_c2_8fc1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2478_c2_8fc1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2478_c2_8fc1]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2491_c11_5d9c]
signal BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2491_c7_8250]
signal t8_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2491_c7_8250]
signal n8_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2491_c7_8250]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2491_c7_8250]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2491_c7_8250]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2491_c7_8250]
signal result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2491_c7_8250]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2494_c11_f758]
signal BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2494_c7_e37a]
signal t8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2494_c7_e37a]
signal n8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2494_c7_e37a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2494_c7_e37a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2494_c7_e37a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2494_c7_e37a]
signal result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2494_c7_e37a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2497_c11_bc34]
signal BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2497_c7_c12d]
signal n8_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2497_c7_c12d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2497_c7_c12d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2497_c7_c12d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2497_c7_c12d]
signal result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2497_c7_c12d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2499_c30_c6da]
signal sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2502_c21_21df]
signal BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_188e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_ram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee
BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_left,
BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_right,
BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output);

-- t8_MUX_uxn_opcodes_h_l2478_c2_8fc1
t8_MUX_uxn_opcodes_h_l2478_c2_8fc1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond,
t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue,
t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse,
t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

-- n8_MUX_uxn_opcodes_h_l2478_c2_8fc1
n8_MUX_uxn_opcodes_h_l2478_c2_8fc1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond,
n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue,
n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse,
n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1
result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1
result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1
result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1
result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1
result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1
result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1
result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c
BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_left,
BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_right,
BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output);

-- t8_MUX_uxn_opcodes_h_l2491_c7_8250
t8_MUX_uxn_opcodes_h_l2491_c7_8250 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2491_c7_8250_cond,
t8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue,
t8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse,
t8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output);

-- n8_MUX_uxn_opcodes_h_l2491_c7_8250
n8_MUX_uxn_opcodes_h_l2491_c7_8250 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2491_c7_8250_cond,
n8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue,
n8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse,
n8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250
result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250
result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250
result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_cond,
result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250
result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758
BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_left,
BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_right,
BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output);

-- t8_MUX_uxn_opcodes_h_l2494_c7_e37a
t8_MUX_uxn_opcodes_h_l2494_c7_e37a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond,
t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue,
t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse,
t8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output);

-- n8_MUX_uxn_opcodes_h_l2494_c7_e37a
n8_MUX_uxn_opcodes_h_l2494_c7_e37a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond,
n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue,
n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse,
n8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a
result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a
result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a
result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34
BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_left,
BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_right,
BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output);

-- n8_MUX_uxn_opcodes_h_l2497_c7_c12d
n8_MUX_uxn_opcodes_h_l2497_c7_c12d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2497_c7_c12d_cond,
n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue,
n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse,
n8_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d
result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d
result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d
result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da
sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_ins,
sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_x,
sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_y,
sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df
BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_left,
BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_right,
BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output,
 t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
 n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output,
 t8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output,
 n8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output,
 t8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output,
 n8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output,
 n8_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output,
 sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2483_c3_e68a : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2488_c3_d5b6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2492_c3_750d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2501_c3_4bce : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2478_l2497_l2491_l2494_DUPLICATE_6f63_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_a0c9_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_84e8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_dcbb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2497_l2494_DUPLICATE_a5e5_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2506_l2474_DUPLICATE_21a7_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2488_c3_d5b6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2488_c3_d5b6;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2483_c3_e68a := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2483_c3_e68a;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2492_c3_750d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2492_c3_750d;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2501_c3_4bce := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2501_c3_4bce;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_a0c9 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_a0c9_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2497_c11_bc34] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_left;
     BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output := BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2502_c21_21df] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_dcbb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_dcbb_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2478_c6_46ee] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_left;
     BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output := BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output := result.is_vram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_84e8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_84e8_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l2499_c30_c6da] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_ins;
     sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_x;
     sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_return_output := sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2497_l2494_DUPLICATE_a5e5 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2497_l2494_DUPLICATE_a5e5_return_output := result.stack_address_sp_offset;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2478_l2497_l2491_l2494_DUPLICATE_6f63 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2478_l2497_l2491_l2494_DUPLICATE_6f63_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2494_c11_f758] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_left;
     BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output := BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2491_c11_5d9c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2478_c6_46ee_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2491_c11_5d9c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2494_c11_f758_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2497_c11_bc34_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2502_c21_21df_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_a0c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_a0c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_a0c9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_dcbb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_dcbb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_dcbb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_84e8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_84e8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2497_l2491_l2494_DUPLICATE_84e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2497_l2494_DUPLICATE_a5e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2497_l2494_DUPLICATE_a5e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2478_l2497_l2491_l2494_DUPLICATE_6f63_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2478_l2497_l2491_l2494_DUPLICATE_6f63_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2478_l2497_l2491_l2494_DUPLICATE_6f63_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2478_l2497_l2491_l2494_DUPLICATE_6f63_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2478_c2_8fc1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2499_c30_c6da_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2497_c7_c12d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2497_c7_c12d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2497_c7_c12d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2497_c7_c12d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_cond;
     n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue;
     n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output := n8_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;

     -- t8_MUX[uxn_opcodes_h_l2494_c7_e37a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond <= VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond;
     t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue;
     t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output := t8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2497_c7_c12d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2497_c7_c12d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2497_c7_c12d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2497_c7_c12d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2494_c7_e37a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2494_c7_e37a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2494_c7_e37a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;

     -- n8_MUX[uxn_opcodes_h_l2494_c7_e37a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_cond;
     n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue;
     n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output := n8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2494_c7_e37a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2494_c7_e37a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;

     -- t8_MUX[uxn_opcodes_h_l2491_c7_8250] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2491_c7_8250_cond <= VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_cond;
     t8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue;
     t8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output := t8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2494_c7_e37a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2491_c7_8250] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;

     -- n8_MUX[uxn_opcodes_h_l2491_c7_8250] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2491_c7_8250_cond <= VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_cond;
     n8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue;
     n8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output := n8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2491_c7_8250] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_return_output := result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2491_c7_8250] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2491_c7_8250] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;

     -- t8_MUX[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond <= VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond;
     t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue;
     t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output := t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2491_c7_8250] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2491_c7_8250_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;
     -- n8_MUX[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond <= VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond;
     n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue;
     n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output := n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2478_c2_8fc1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2506_l2474_DUPLICATE_21a7 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2506_l2474_DUPLICATE_21a7_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_188e(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2478_c2_8fc1_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2506_l2474_DUPLICATE_21a7_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2506_l2474_DUPLICATE_21a7_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
