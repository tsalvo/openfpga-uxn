-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity dup2_0CLK_e4095020 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup2_0CLK_e4095020;
architecture arch of dup2_0CLK_e4095020 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2790_c6_b17a]
signal BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2790_c2_065c]
signal t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2790_c2_065c]
signal t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2790_c2_065c]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2790_c2_065c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2790_c2_065c]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2790_c2_065c]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2790_c2_065c]
signal result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2790_c2_065c]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2790_c2_065c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2790_c2_065c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2790_c2_065c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2803_c11_086a]
signal BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2803_c7_f28d]
signal t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2803_c7_f28d]
signal t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2803_c7_f28d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2803_c7_f28d]
signal result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2803_c7_f28d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2803_c7_f28d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2803_c7_f28d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2806_c11_cbf9]
signal BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2806_c7_b3e8]
signal t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2806_c7_b3e8]
signal t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2806_c7_b3e8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2806_c7_b3e8]
signal result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2806_c7_b3e8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2806_c7_b3e8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2806_c7_b3e8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2808_c30_1948]
signal sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2813_c11_19c5]
signal BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2813_c7_18e3]
signal t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2813_c7_18e3]
signal result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2813_c7_18e3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2813_c7_18e3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2813_c7_18e3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2819_c11_c4f9]
signal BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2819_c7_89c9]
signal result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2819_c7_89c9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2819_c7_89c9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2823_c11_59d4]
signal BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2823_c7_befb]
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2823_c7_befb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2823_c7_befb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_return_output : unsigned(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a
BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_left,
BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_right,
BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2790_c2_065c
t16_low_MUX_uxn_opcodes_h_l2790_c2_065c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_cond,
t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue,
t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse,
t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2790_c2_065c
t16_high_MUX_uxn_opcodes_h_l2790_c2_065c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_cond,
t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue,
t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse,
t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c
result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c
result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c
result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c
result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c
result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c
result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a
BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_left,
BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_right,
BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d
t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_cond,
t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue,
t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse,
t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d
t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_cond,
t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue,
t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse,
t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d
result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d
result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d
result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9
BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_left,
BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_right,
BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8
t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond,
t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue,
t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse,
t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8
t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond,
t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue,
t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse,
t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8
result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8
result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8
result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2808_c30_1948
sp_relative_shift_uxn_opcodes_h_l2808_c30_1948 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_ins,
sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_x,
sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_y,
sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5
BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_left,
BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_right,
BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3
t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_cond,
t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue,
t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse,
t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3
result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3
result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9
BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_left,
BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_right,
BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9
result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9
result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_left,
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_right,
BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_cond,
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output,
 t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
 t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output,
 t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output,
 t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output,
 t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output,
 t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output,
 sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_return_output,
 t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2795_c3_9cb9 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2800_c3_950d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2804_c3_e88d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2810_c3_f784 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2815_c3_9f73 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2816_c3_952a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2820_c3_2ad3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2824_c3_6c9b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2823_c7_befb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_87be_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2803_l2806_DUPLICATE_941f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2803_l2813_DUPLICATE_621c_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2823_l2819_l2813_l2806_l2803_DUPLICATE_49e7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2786_l2829_DUPLICATE_62cd_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2816_c3_952a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2816_c3_952a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_right := to_unsigned(5, 3);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2804_c3_e88d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2804_c3_e88d;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_right := to_unsigned(4, 3);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2815_c3_9f73 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2815_c3_9f73;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2795_c3_9cb9 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2795_c3_9cb9;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2820_c3_2ad3 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2820_c3_2ad3;
     VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2810_c3_f784 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2810_c3_f784;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_y := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2824_c3_6c9b := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2824_c3_6c9b;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2800_c3_950d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2800_c3_950d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse := t16_low;
     -- BIN_OP_EQ[uxn_opcodes_h_l2819_c11_c4f9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2790_c2_065c_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2813_c11_19c5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2790_c2_065c_return_output := result.is_pc_updated;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2790_c2_065c_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2803_l2806_DUPLICATE_941f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2803_l2806_DUPLICATE_941f_return_output := result.is_stack_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2823_c7_befb] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2823_c7_befb_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2790_c6_b17a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2823_c11_59d4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2806_c11_cbf9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2790_c2_065c_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2823_l2819_l2813_l2806_l2803_DUPLICATE_49e7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2823_l2819_l2813_l2806_l2803_DUPLICATE_49e7_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2803_l2813_DUPLICATE_621c LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2803_l2813_DUPLICATE_621c_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2803_c11_086a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2808_c30_1948] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_ins;
     sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_x;
     sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_return_output := sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_87be LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_87be_return_output := result.u8_value;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2790_c6_b17a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2803_c11_086a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2806_c11_cbf9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2813_c11_19c5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2819_c11_c4f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2823_c11_59d4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2803_l2813_DUPLICATE_621c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2803_l2813_DUPLICATE_621c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2823_l2819_l2813_l2806_l2803_DUPLICATE_49e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2823_l2819_l2813_l2806_l2803_DUPLICATE_49e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2823_l2819_l2813_l2806_l2803_DUPLICATE_49e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2823_l2819_l2813_l2806_l2803_DUPLICATE_49e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2823_l2819_l2813_l2806_l2803_DUPLICATE_49e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2803_l2806_DUPLICATE_941f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2803_l2806_DUPLICATE_941f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_87be_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_87be_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2803_l2823_l2790_DUPLICATE_87be_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2790_c2_065c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2790_c2_065c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2790_c2_065c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2790_c2_065c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2823_c7_befb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2808_c30_1948_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2813_c7_18e3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2806_c7_b3e8] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond;
     t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output := t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2823_c7_befb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2813_c7_18e3] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_cond;
     t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output := t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2823_c7_befb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2823_c7_befb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_return_output := result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2806_c7_b3e8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2823_c7_befb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2823_c7_befb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2823_c7_befb_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2803_c7_f28d] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_cond;
     t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output := t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2806_c7_b3e8] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond;
     t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output := t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2819_c7_89c9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2819_c7_89c9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2806_c7_b3e8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2803_c7_f28d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2819_c7_89c9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2819_c7_89c9_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;
     -- t16_low_MUX[uxn_opcodes_h_l2803_c7_f28d] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_cond;
     t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output := t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_cond;
     t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_return_output := t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2803_c7_f28d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2813_c7_18e3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2813_c7_18e3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2813_c7_18e3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2813_c7_18e3_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2806_c7_b3e8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2806_c7_b3e8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2806_c7_b3e8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_cond;
     t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_return_output := t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2806_c7_b3e8_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2803_c7_f28d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2803_c7_f28d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2803_c7_f28d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2803_c7_f28d_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2790_c2_065c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2786_l2829_DUPLICATE_62cd LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2786_l2829_DUPLICATE_62cd_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2790_c2_065c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2790_c2_065c_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2786_l2829_DUPLICATE_62cd_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l2786_l2829_DUPLICATE_62cd_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
