-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 41
entity jmp2_0CLK_0b1ee796 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jmp2_0CLK_0b1ee796;
architecture arch of jmp2_0CLK_0b1ee796 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l612_c6_8086]
signal BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l612_c1_b492]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l612_c2_1ccf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l612_c2_1ccf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l612_c2_1ccf]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l612_c2_1ccf]
signal result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l612_c2_1ccf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l612_c2_1ccf]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l612_c2_1ccf]
signal t16_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l613_c3_bf7c[uxn_opcodes_h_l613_c3_bf7c]
signal printf_uxn_opcodes_h_l613_c3_bf7c_uxn_opcodes_h_l613_c3_bf7c_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l617_c11_d1d6]
signal BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l617_c7_a337]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l617_c7_a337]
signal result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l617_c7_a337]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l617_c7_a337]
signal result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l617_c7_a337]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l617_c7_a337]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l617_c7_a337]
signal t16_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l620_c11_45dc]
signal BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l620_c7_f2b1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l620_c7_f2b1]
signal result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l620_c7_f2b1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l620_c7_f2b1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l620_c7_f2b1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l620_c7_f2b1]
signal t16_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l622_c3_8f90]
signal CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l624_c11_e5bf]
signal BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l624_c7_04ff]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l624_c7_04ff]
signal result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l624_c7_04ff]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l624_c7_04ff]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l624_c7_04ff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l624_c7_04ff]
signal t16_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l625_c3_a865]
signal BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l627_c30_d9bc]
signal sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l631_c11_5d87]
signal BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l631_c7_2587]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l631_c7_2587]
signal result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l631_c7_2587]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_5d97( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.u16_value := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_pc_updated := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086
BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_left,
BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_right,
BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf
result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf
result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf
result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_cond,
result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf
result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf
result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output);

-- t16_MUX_uxn_opcodes_h_l612_c2_1ccf
t16_MUX_uxn_opcodes_h_l612_c2_1ccf : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l612_c2_1ccf_cond,
t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue,
t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse,
t16_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output);

-- printf_uxn_opcodes_h_l613_c3_bf7c_uxn_opcodes_h_l613_c3_bf7c
printf_uxn_opcodes_h_l613_c3_bf7c_uxn_opcodes_h_l613_c3_bf7c : entity work.printf_uxn_opcodes_h_l613_c3_bf7c_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l613_c3_bf7c_uxn_opcodes_h_l613_c3_bf7c_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6
BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_left,
BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_right,
BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337
result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337
result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337
result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_cond,
result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337
result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337
result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_return_output);

-- t16_MUX_uxn_opcodes_h_l617_c7_a337
t16_MUX_uxn_opcodes_h_l617_c7_a337 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l617_c7_a337_cond,
t16_MUX_uxn_opcodes_h_l617_c7_a337_iftrue,
t16_MUX_uxn_opcodes_h_l617_c7_a337_iffalse,
t16_MUX_uxn_opcodes_h_l617_c7_a337_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc
BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_left,
BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_right,
BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1
result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1
result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_cond,
result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1
result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1
result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1
result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output);

-- t16_MUX_uxn_opcodes_h_l620_c7_f2b1
t16_MUX_uxn_opcodes_h_l620_c7_f2b1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l620_c7_f2b1_cond,
t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue,
t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse,
t16_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output);

-- CONST_SL_8_uxn_opcodes_h_l622_c3_8f90
CONST_SL_8_uxn_opcodes_h_l622_c3_8f90 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_x,
CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf
BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_left,
BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_right,
BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff
result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff
result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_cond,
result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff
result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff
result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff
result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_return_output);

-- t16_MUX_uxn_opcodes_h_l624_c7_04ff
t16_MUX_uxn_opcodes_h_l624_c7_04ff : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l624_c7_04ff_cond,
t16_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue,
t16_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse,
t16_MUX_uxn_opcodes_h_l624_c7_04ff_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l625_c3_a865
BIN_OP_OR_uxn_opcodes_h_l625_c3_a865 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_left,
BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_right,
BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_return_output);

-- sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc
sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_ins,
sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_x,
sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_y,
sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87
BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_left,
BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_right,
BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587
result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587
result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587
result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
 t16_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_return_output,
 t16_MUX_uxn_opcodes_h_l617_c7_a337_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output,
 t16_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output,
 CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_return_output,
 t16_MUX_uxn_opcodes_h_l624_c7_04ff_return_output,
 BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_return_output,
 sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l614_c3_57a9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l613_c3_bf7c_uxn_opcodes_h_l613_c3_bf7c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l618_c3_bb81 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l617_c7_a337_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_return_output : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_bec5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_59b4_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_1572_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_88e1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l617_l631_l620_l624_DUPLICATE_6459_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l625_l621_DUPLICATE_8092_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5d97_uxn_opcodes_h_l608_l637_DUPLICATE_0554_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l618_c3_bb81 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l618_c3_bb81;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l614_c3_57a9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l614_c3_57a9;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l617_c11_d1d6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_left;
     BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output := BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l612_c6_8086] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_left;
     BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output := BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l620_c11_45dc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_left;
     BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output := BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_88e1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_88e1_return_output := result.is_pc_updated;

     -- sp_relative_shift[uxn_opcodes_h_l627_c30_d9bc] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_ins;
     sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_x <= VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_x;
     sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_y <= VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_return_output := sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l617_l631_l620_l624_DUPLICATE_6459 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l617_l631_l620_l624_DUPLICATE_6459_return_output := result.is_opc_done;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l617_c7_a337] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l617_c7_a337_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l631_c11_5d87] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_left;
     BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_return_output := BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_1572 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_1572_return_output := result.sp_relative_shift;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l625_l621_DUPLICATE_8092 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l625_l621_DUPLICATE_8092_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l624_c11_e5bf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_left;
     BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output := BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_bec5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_bec5_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_59b4 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_59b4_return_output := result.u16_value;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l612_c6_8086_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l617_c11_d1d6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l620_c11_45dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l624_c11_e5bf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l631_c11_5d87_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l625_l621_DUPLICATE_8092_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l625_l621_DUPLICATE_8092_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_1572_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_1572_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_1572_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_1572_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_59b4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_59b4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_59b4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l617_l620_l612_l624_DUPLICATE_59b4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l617_l631_l620_l624_DUPLICATE_6459_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l617_l631_l620_l624_DUPLICATE_6459_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l617_l631_l620_l624_DUPLICATE_6459_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l617_l631_l620_l624_DUPLICATE_6459_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_88e1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_88e1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_88e1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_88e1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_bec5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_bec5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_bec5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l617_l631_l620_l612_DUPLICATE_bec5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l617_c7_a337_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l627_c30_d9bc_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l631_c7_2587] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l622_c3_8f90] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_x <= VAR_CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_return_output := CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l612_c1_b492] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l617_c7_a337] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l624_c7_04ff] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l625_c3_a865] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_left;
     BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_return_output := BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l631_c7_2587] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l631_c7_2587] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_return_output;

     -- Submodule level 2
     VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l625_c3_a865_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l622_c3_8f90_return_output;
     VAR_printf_uxn_opcodes_h_l613_c3_bf7c_uxn_opcodes_h_l613_c3_bf7c_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l612_c1_b492_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l631_c7_2587_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l631_c7_2587_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l631_c7_2587_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l617_c7_a337_return_output;
     -- printf_uxn_opcodes_h_l613_c3_bf7c[uxn_opcodes_h_l613_c3_bf7c] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l613_c3_bf7c_uxn_opcodes_h_l613_c3_bf7c_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l613_c3_bf7c_uxn_opcodes_h_l613_c3_bf7c_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t16_MUX[uxn_opcodes_h_l624_c7_04ff] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l624_c7_04ff_cond <= VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_cond;
     t16_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue;
     t16_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_return_output := t16_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l624_c7_04ff] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_cond;
     result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_return_output := result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l624_c7_04ff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l624_c7_04ff] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l624_c7_04ff] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l612_c2_1ccf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l620_c7_f2b1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse := VAR_t16_MUX_uxn_opcodes_h_l624_c7_04ff_return_output;
     -- t16_MUX[uxn_opcodes_h_l620_c7_f2b1] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l620_c7_f2b1_cond <= VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_cond;
     t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue;
     t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output := t16_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l620_c7_f2b1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l620_c7_f2b1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l620_c7_f2b1] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_cond;
     result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output := result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l617_c7_a337] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l620_c7_f2b1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_iffalse := VAR_t16_MUX_uxn_opcodes_h_l620_c7_f2b1_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l617_c7_a337] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l617_c7_a337] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l612_c2_1ccf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output;

     -- t16_MUX[uxn_opcodes_h_l617_c7_a337] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l617_c7_a337_cond <= VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_cond;
     t16_MUX_uxn_opcodes_h_l617_c7_a337_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_iftrue;
     t16_MUX_uxn_opcodes_h_l617_c7_a337_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_return_output := t16_MUX_uxn_opcodes_h_l617_c7_a337_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l617_c7_a337] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_cond;
     result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_return_output := result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l617_c7_a337] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l617_c7_a337_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l617_c7_a337_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l617_c7_a337_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l617_c7_a337_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse := VAR_t16_MUX_uxn_opcodes_h_l617_c7_a337_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l612_c2_1ccf] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output;

     -- t16_MUX[uxn_opcodes_h_l612_c2_1ccf] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l612_c2_1ccf_cond <= VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_cond;
     t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue;
     t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output := t16_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l612_c2_1ccf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l612_c2_1ccf] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_cond;
     result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output := result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l612_c2_1ccf] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output;

     -- Submodule level 6
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5d97_uxn_opcodes_h_l608_l637_DUPLICATE_0554 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5d97_uxn_opcodes_h_l608_l637_DUPLICATE_0554_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5d97(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l612_c2_1ccf_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5d97_uxn_opcodes_h_l608_l637_DUPLICATE_0554_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5d97_uxn_opcodes_h_l608_l637_DUPLICATE_0554_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
