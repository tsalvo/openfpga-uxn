-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity jcn2_0CLK_db1e6fcb is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jcn2_0CLK_db1e6fcb;
architecture arch of jcn2_0CLK_db1e6fcb is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l684_c6_e2bf]
signal BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l684_c2_d22f]
signal n8_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l684_c2_d22f]
signal t16_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l684_c2_d22f]
signal result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l684_c2_d22f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l684_c2_d22f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l684_c2_d22f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l684_c2_d22f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l691_c11_2f0c]
signal BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l691_c7_3b7a]
signal n8_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l691_c7_3b7a]
signal t16_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l691_c7_3b7a]
signal result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l691_c7_3b7a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l691_c7_3b7a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l691_c7_3b7a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l691_c7_3b7a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l694_c11_2ec8]
signal BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l694_c7_7342]
signal n8_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l694_c7_7342]
signal t16_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l694_c7_7342]
signal result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l694_c7_7342]
signal result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l694_c7_7342]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l694_c7_7342]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l694_c7_7342]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(3 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l696_c3_21e5]
signal CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l699_c11_2c7d]
signal BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l699_c7_c9bd]
signal n8_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l699_c7_c9bd]
signal t16_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l699_c7_c9bd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l699_c7_c9bd]
signal result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l699_c7_c9bd]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l699_c7_c9bd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l700_c3_2852]
signal BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l702_c11_15a2]
signal BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l702_c7_4202]
signal n8_MUX_uxn_opcodes_h_l702_c7_4202_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l702_c7_4202_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l702_c7_4202_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l702_c7_4202_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l702_c7_4202]
signal result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l702_c7_4202]
signal result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l702_c7_4202]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l702_c7_4202]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l705_c30_b6e3]
signal sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l706_c26_a7e1]
signal BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l706_c26_a9b9]
signal MUX_uxn_opcodes_h_l706_c26_a9b9_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l706_c26_a9b9_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l706_c26_a9b9_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l706_c26_a9b9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l707_c22_42f0]
signal BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l707_c22_11f7]
signal MUX_uxn_opcodes_h_l707_c22_11f7_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l707_c22_11f7_iftrue : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l707_c22_11f7_iffalse : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l707_c22_11f7_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l709_c11_f23e]
signal BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l709_c7_68b5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l709_c7_68b5]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l709_c7_68b5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_return_output : signed(3 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_6e0b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.is_pc_updated := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf
BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_left,
BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_right,
BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output);

-- n8_MUX_uxn_opcodes_h_l684_c2_d22f
n8_MUX_uxn_opcodes_h_l684_c2_d22f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l684_c2_d22f_cond,
n8_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue,
n8_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse,
n8_MUX_uxn_opcodes_h_l684_c2_d22f_return_output);

-- t16_MUX_uxn_opcodes_h_l684_c2_d22f
t16_MUX_uxn_opcodes_h_l684_c2_d22f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l684_c2_d22f_cond,
t16_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue,
t16_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse,
t16_MUX_uxn_opcodes_h_l684_c2_d22f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f
result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_cond,
result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f
result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f
result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f
result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c
BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_left,
BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_right,
BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output);

-- n8_MUX_uxn_opcodes_h_l691_c7_3b7a
n8_MUX_uxn_opcodes_h_l691_c7_3b7a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l691_c7_3b7a_cond,
n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue,
n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse,
n8_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output);

-- t16_MUX_uxn_opcodes_h_l691_c7_3b7a
t16_MUX_uxn_opcodes_h_l691_c7_3b7a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l691_c7_3b7a_cond,
t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue,
t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse,
t16_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a
result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_cond,
result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a
result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a
result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a
result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8
BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_left,
BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_right,
BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output);

-- n8_MUX_uxn_opcodes_h_l694_c7_7342
n8_MUX_uxn_opcodes_h_l694_c7_7342 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l694_c7_7342_cond,
n8_MUX_uxn_opcodes_h_l694_c7_7342_iftrue,
n8_MUX_uxn_opcodes_h_l694_c7_7342_iffalse,
n8_MUX_uxn_opcodes_h_l694_c7_7342_return_output);

-- t16_MUX_uxn_opcodes_h_l694_c7_7342
t16_MUX_uxn_opcodes_h_l694_c7_7342 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l694_c7_7342_cond,
t16_MUX_uxn_opcodes_h_l694_c7_7342_iftrue,
t16_MUX_uxn_opcodes_h_l694_c7_7342_iffalse,
t16_MUX_uxn_opcodes_h_l694_c7_7342_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342
result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_cond,
result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342
result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342
result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342
result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_return_output);

-- CONST_SL_8_uxn_opcodes_h_l696_c3_21e5
CONST_SL_8_uxn_opcodes_h_l696_c3_21e5 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_x,
CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d
BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_left,
BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_right,
BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output);

-- n8_MUX_uxn_opcodes_h_l699_c7_c9bd
n8_MUX_uxn_opcodes_h_l699_c7_c9bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l699_c7_c9bd_cond,
n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue,
n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse,
n8_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output);

-- t16_MUX_uxn_opcodes_h_l699_c7_c9bd
t16_MUX_uxn_opcodes_h_l699_c7_c9bd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l699_c7_c9bd_cond,
t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue,
t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse,
t16_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd
result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd
result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_cond,
result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd
result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd
result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l700_c3_2852
BIN_OP_OR_uxn_opcodes_h_l700_c3_2852 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_left,
BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_right,
BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2
BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_left,
BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_right,
BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_return_output);

-- n8_MUX_uxn_opcodes_h_l702_c7_4202
n8_MUX_uxn_opcodes_h_l702_c7_4202 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l702_c7_4202_cond,
n8_MUX_uxn_opcodes_h_l702_c7_4202_iftrue,
n8_MUX_uxn_opcodes_h_l702_c7_4202_iffalse,
n8_MUX_uxn_opcodes_h_l702_c7_4202_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202
result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202
result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_cond,
result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202
result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202
result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_return_output);

-- sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3
sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_ins,
sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_x,
sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_y,
sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1
BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_left,
BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_right,
BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_return_output);

-- MUX_uxn_opcodes_h_l706_c26_a9b9
MUX_uxn_opcodes_h_l706_c26_a9b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l706_c26_a9b9_cond,
MUX_uxn_opcodes_h_l706_c26_a9b9_iftrue,
MUX_uxn_opcodes_h_l706_c26_a9b9_iffalse,
MUX_uxn_opcodes_h_l706_c26_a9b9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0
BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_left,
BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_right,
BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_return_output);

-- MUX_uxn_opcodes_h_l707_c22_11f7
MUX_uxn_opcodes_h_l707_c22_11f7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l707_c22_11f7_cond,
MUX_uxn_opcodes_h_l707_c22_11f7_iftrue,
MUX_uxn_opcodes_h_l707_c22_11f7_iffalse,
MUX_uxn_opcodes_h_l707_c22_11f7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e
BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_left,
BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_right,
BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5
result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5
result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5
result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output,
 n8_MUX_uxn_opcodes_h_l684_c2_d22f_return_output,
 t16_MUX_uxn_opcodes_h_l684_c2_d22f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output,
 n8_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output,
 t16_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output,
 n8_MUX_uxn_opcodes_h_l694_c7_7342_return_output,
 t16_MUX_uxn_opcodes_h_l694_c7_7342_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_return_output,
 CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output,
 n8_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output,
 t16_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output,
 BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_return_output,
 n8_MUX_uxn_opcodes_h_l702_c7_4202_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_return_output,
 sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_return_output,
 MUX_uxn_opcodes_h_l706_c26_a9b9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_return_output,
 MUX_uxn_opcodes_h_l707_c22_11f7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l688_c3_1c43 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l692_c3_de5e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l697_c3_d7ea : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l694_c7_7342_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l707_c22_11f7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l707_c22_11f7_iftrue : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l707_c22_11f7_iffalse : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l707_c22_11f7_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l710_c3_cd1d : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l702_l699_l694_l691_l684_DUPLICATE_ce6b_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_c317_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_b078_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l702_l699_l694_l691_l709_DUPLICATE_5e32_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l700_l695_DUPLICATE_950a_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6e0b_uxn_opcodes_h_l679_l715_DUPLICATE_6fb0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_opcodes_h_l707_c22_11f7_iftrue := resize(to_unsigned(0, 1), 16);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_y := resize(to_signed(-3, 3), 4);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l710_c3_cd1d := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l710_c3_cd1d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_right := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_iffalse := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l688_c3_1c43 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l688_c3_1c43;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l697_c3_d7ea := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l697_c3_d7ea;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l692_c3_de5e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l692_c3_de5e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_left := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_left := t16;
     VAR_MUX_uxn_opcodes_h_l707_c22_11f7_iffalse := t16;
     VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse := t16;
     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l700_l695_DUPLICATE_950a LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l700_l695_DUPLICATE_950a_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l694_c11_2ec8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_left;
     BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output := BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l702_l699_l694_l691_l684_DUPLICATE_ce6b LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l702_l699_l694_l691_l684_DUPLICATE_ce6b_return_output := result.u16_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l694_c7_7342] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l694_c7_7342_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l691_c11_2f0c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_left;
     BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output := BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_c317 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_c317_return_output := result.is_pc_updated;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_b078 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_b078_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l706_c26_a7e1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_left;
     BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_return_output := BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l702_c11_15a2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_left;
     BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_return_output := BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l709_c11_f23e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_left;
     BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_return_output := BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l702_l699_l694_l691_l709_DUPLICATE_5e32 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l702_l699_l694_l691_l709_DUPLICATE_5e32_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l705_c30_b6e3] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_ins;
     sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_x <= VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_x;
     sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_y <= VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_return_output := sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l707_c22_42f0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_left;
     BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_return_output := BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l684_c6_e2bf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_left;
     BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output := BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l699_c11_2c7d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_left;
     BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output := BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l684_c6_e2bf_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l691_c11_2f0c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l694_c11_2ec8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l699_c11_2c7d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l702_c11_15a2_return_output;
     VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l706_c26_a7e1_return_output;
     VAR_MUX_uxn_opcodes_h_l707_c22_11f7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l707_c22_42f0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l709_c11_f23e_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l700_l695_DUPLICATE_950a_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l700_l695_DUPLICATE_950a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_b078_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_b078_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_b078_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_b078_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_b078_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l702_l699_l694_l691_l684_DUPLICATE_ce6b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l702_l699_l694_l691_l684_DUPLICATE_ce6b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l702_l699_l694_l691_l684_DUPLICATE_ce6b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l702_l699_l694_l691_l684_DUPLICATE_ce6b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l702_l699_l694_l691_l684_DUPLICATE_ce6b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l702_l699_l694_l691_l709_DUPLICATE_5e32_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l702_l699_l694_l691_l709_DUPLICATE_5e32_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l702_l699_l694_l691_l709_DUPLICATE_5e32_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l702_l699_l694_l691_l709_DUPLICATE_5e32_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l702_l699_l694_l691_l709_DUPLICATE_5e32_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_c317_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_c317_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_c317_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_c317_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l699_l694_l691_l684_l709_DUPLICATE_c317_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l694_c7_7342_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l705_c30_b6e3_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l709_c7_68b5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l696_c3_21e5] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_x <= VAR_CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_return_output := CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_return_output;

     -- MUX[uxn_opcodes_h_l706_c26_a9b9] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l706_c26_a9b9_cond <= VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_cond;
     MUX_uxn_opcodes_h_l706_c26_a9b9_iftrue <= VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_iftrue;
     MUX_uxn_opcodes_h_l706_c26_a9b9_iffalse <= VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_return_output := MUX_uxn_opcodes_h_l706_c26_a9b9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l709_c7_68b5] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l700_c3_2852] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_left;
     BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_return_output := BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l709_c7_68b5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l694_c7_7342] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_return_output;

     -- MUX[uxn_opcodes_h_l707_c22_11f7] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l707_c22_11f7_cond <= VAR_MUX_uxn_opcodes_h_l707_c22_11f7_cond;
     MUX_uxn_opcodes_h_l707_c22_11f7_iftrue <= VAR_MUX_uxn_opcodes_h_l707_c22_11f7_iftrue;
     MUX_uxn_opcodes_h_l707_c22_11f7_iffalse <= VAR_MUX_uxn_opcodes_h_l707_c22_11f7_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l707_c22_11f7_return_output := MUX_uxn_opcodes_h_l707_c22_11f7_return_output;

     -- n8_MUX[uxn_opcodes_h_l702_c7_4202] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l702_c7_4202_cond <= VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_cond;
     n8_MUX_uxn_opcodes_h_l702_c7_4202_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_iftrue;
     n8_MUX_uxn_opcodes_h_l702_c7_4202_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_return_output := n8_MUX_uxn_opcodes_h_l702_c7_4202_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l700_c3_2852_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l696_c3_21e5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iftrue := VAR_MUX_uxn_opcodes_h_l706_c26_a9b9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iftrue := VAR_MUX_uxn_opcodes_h_l707_c22_11f7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l702_c7_4202_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l709_c7_68b5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l709_c7_68b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l709_c7_68b5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l694_c7_7342_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l702_c7_4202] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_cond;
     result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_return_output := result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l691_c7_3b7a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l702_c7_4202] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_return_output;

     -- n8_MUX[uxn_opcodes_h_l699_c7_c9bd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l699_c7_c9bd_cond <= VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_cond;
     n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue;
     n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output := n8_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l702_c7_4202] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_return_output;

     -- t16_MUX[uxn_opcodes_h_l699_c7_c9bd] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l699_c7_c9bd_cond <= VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_cond;
     t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue;
     t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output := t16_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l702_c7_4202] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_iffalse := VAR_n8_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l702_c7_4202_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l702_c7_4202_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l702_c7_4202_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l702_c7_4202_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_iffalse := VAR_t16_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;
     -- n8_MUX[uxn_opcodes_h_l694_c7_7342] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l694_c7_7342_cond <= VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_cond;
     n8_MUX_uxn_opcodes_h_l694_c7_7342_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_iftrue;
     n8_MUX_uxn_opcodes_h_l694_c7_7342_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_return_output := n8_MUX_uxn_opcodes_h_l694_c7_7342_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l699_c7_c9bd] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_cond;
     result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output := result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l699_c7_c9bd] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l699_c7_c9bd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l699_c7_c9bd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;

     -- t16_MUX[uxn_opcodes_h_l694_c7_7342] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l694_c7_7342_cond <= VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_cond;
     t16_MUX_uxn_opcodes_h_l694_c7_7342_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_iftrue;
     t16_MUX_uxn_opcodes_h_l694_c7_7342_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_return_output := t16_MUX_uxn_opcodes_h_l694_c7_7342_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l684_c2_d22f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l694_c7_7342_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l699_c7_c9bd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse := VAR_t16_MUX_uxn_opcodes_h_l694_c7_7342_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l694_c7_7342] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_return_output;

     -- n8_MUX[uxn_opcodes_h_l691_c7_3b7a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l691_c7_3b7a_cond <= VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_cond;
     n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue;
     n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output := n8_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l694_c7_7342] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l694_c7_7342] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l694_c7_7342] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_cond;
     result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_return_output := result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_return_output;

     -- t16_MUX[uxn_opcodes_h_l691_c7_3b7a] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l691_c7_3b7a_cond <= VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_cond;
     t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue;
     t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output := t16_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l694_c7_7342_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l694_c7_7342_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l694_c7_7342_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l694_c7_7342_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse := VAR_t16_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l691_c7_3b7a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l691_c7_3b7a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;

     -- n8_MUX[uxn_opcodes_h_l684_c2_d22f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l684_c2_d22f_cond <= VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_cond;
     n8_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue;
     n8_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_return_output := n8_MUX_uxn_opcodes_h_l684_c2_d22f_return_output;

     -- t16_MUX[uxn_opcodes_h_l684_c2_d22f] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l684_c2_d22f_cond <= VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_cond;
     t16_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue;
     t16_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_return_output := t16_MUX_uxn_opcodes_h_l684_c2_d22f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l691_c7_3b7a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output := result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l691_c7_3b7a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l684_c2_d22f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l691_c7_3b7a_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l684_c2_d22f_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l684_c2_d22f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l684_c2_d22f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l684_c2_d22f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_return_output := result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l684_c2_d22f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_6e0b_uxn_opcodes_h_l679_l715_DUPLICATE_6fb0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6e0b_uxn_opcodes_h_l679_l715_DUPLICATE_6fb0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_6e0b(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l684_c2_d22f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l684_c2_d22f_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l684_c2_d22f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l684_c2_d22f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l684_c2_d22f_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6e0b_uxn_opcodes_h_l679_l715_DUPLICATE_6fb0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6e0b_uxn_opcodes_h_l679_l715_DUPLICATE_6fb0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
