-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity eor_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_bacf6a1d;
architecture arch of eor_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1035_c6_f247]
signal BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1035_c1_8e35]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1035_c2_df05]
signal t8_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1035_c2_df05]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1035_c2_df05]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1035_c2_df05]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1035_c2_df05]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1035_c2_df05]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1035_c2_df05]
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1035_c2_df05]
signal n8_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1036_c3_dc0e[uxn_opcodes_h_l1036_c3_dc0e]
signal printf_uxn_opcodes_h_l1036_c3_dc0e_uxn_opcodes_h_l1036_c3_dc0e_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1040_c11_2db6]
signal BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1040_c7_fdab]
signal t8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1040_c7_fdab]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1040_c7_fdab]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1040_c7_fdab]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1040_c7_fdab]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1040_c7_fdab]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1040_c7_fdab]
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1040_c7_fdab]
signal n8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1043_c11_fa4a]
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1043_c7_f340]
signal t8_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1043_c7_f340]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1043_c7_f340]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1043_c7_f340]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1043_c7_f340]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1043_c7_f340]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1043_c7_f340]
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1043_c7_f340]
signal n8_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1046_c11_fe55]
signal BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1046_c7_55cd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1046_c7_55cd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1046_c7_55cd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1046_c7_55cd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1046_c7_55cd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1046_c7_55cd]
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1046_c7_55cd]
signal n8_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1049_c30_eb5b]
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1052_c21_cf1e]
signal BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1054_c11_0275]
signal BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1054_c7_5d8c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1054_c7_5d8c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1054_c7_5d8c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8c29( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_left,
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_right,
BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_return_output);

-- t8_MUX_uxn_opcodes_h_l1035_c2_df05
t8_MUX_uxn_opcodes_h_l1035_c2_df05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1035_c2_df05_cond,
t8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue,
t8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse,
t8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_cond,
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_return_output);

-- n8_MUX_uxn_opcodes_h_l1035_c2_df05
n8_MUX_uxn_opcodes_h_l1035_c2_df05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1035_c2_df05_cond,
n8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue,
n8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse,
n8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output);

-- printf_uxn_opcodes_h_l1036_c3_dc0e_uxn_opcodes_h_l1036_c3_dc0e
printf_uxn_opcodes_h_l1036_c3_dc0e_uxn_opcodes_h_l1036_c3_dc0e : entity work.printf_uxn_opcodes_h_l1036_c3_dc0e_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1036_c3_dc0e_uxn_opcodes_h_l1036_c3_dc0e_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_left,
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_right,
BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output);

-- t8_MUX_uxn_opcodes_h_l1040_c7_fdab
t8_MUX_uxn_opcodes_h_l1040_c7_fdab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond,
t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue,
t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse,
t8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_cond,
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output);

-- n8_MUX_uxn_opcodes_h_l1040_c7_fdab
n8_MUX_uxn_opcodes_h_l1040_c7_fdab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond,
n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue,
n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse,
n8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_left,
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_right,
BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output);

-- t8_MUX_uxn_opcodes_h_l1043_c7_f340
t8_MUX_uxn_opcodes_h_l1043_c7_f340 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1043_c7_f340_cond,
t8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue,
t8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse,
t8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_cond,
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_return_output);

-- n8_MUX_uxn_opcodes_h_l1043_c7_f340
n8_MUX_uxn_opcodes_h_l1043_c7_f340 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1043_c7_f340_cond,
n8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue,
n8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse,
n8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_left,
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_right,
BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_cond,
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output);

-- n8_MUX_uxn_opcodes_h_l1046_c7_55cd
n8_MUX_uxn_opcodes_h_l1046_c7_55cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1046_c7_55cd_cond,
n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue,
n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse,
n8_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b
sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_ins,
sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_x,
sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_y,
sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_left,
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_right,
BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_left,
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_right,
BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_return_output,
 t8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
 n8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output,
 t8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output,
 n8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output,
 t8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_return_output,
 n8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output,
 n8_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output,
 sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_b91d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1036_c3_dc0e_uxn_opcodes_h_l1036_c3_dc0e_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1041_c3_c613 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_d1b3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_fe89_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3546_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_0685_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_6504_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_ce39_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_9757_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1060_l1031_DUPLICATE_d824_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_d1b3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1051_c3_d1b3;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_b91d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1037_c3_b91d;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_right := to_unsigned(4, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1041_c3_c613 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1041_c3_c613;
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse := t8;
     -- BIN_OP_XOR[uxn_opcodes_h_l1052_c21_cf1e] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_left;
     BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_return_output := BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3546 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3546_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_0685 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_0685_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_6504 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_6504_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_ce39 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_ce39_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1040_c11_2db6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_fe89 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_fe89_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1054_c11_0275] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_left;
     BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_return_output := BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1049_c30_eb5b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_ins;
     sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_x;
     sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_return_output := sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1043_c11_fa4a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_9757 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_9757_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1035_c6_f247] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_left;
     BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output := BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1046_c11_fe55] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_left;
     BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output := BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1035_c6_f247_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1040_c11_2db6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1043_c11_fa4a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1046_c11_fe55_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1054_c11_0275_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1052_c21_cf1e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_0685_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_0685_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_0685_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_0685_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_ce39_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_ce39_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_ce39_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1054_l1043_l1046_l1040_DUPLICATE_ce39_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_fe89_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_fe89_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_fe89_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_fe89_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3546_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3546_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3546_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1054_l1043_l1035_l1040_DUPLICATE_3546_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_9757_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1043_l1046_DUPLICATE_9757_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_6504_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_6504_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_6504_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1043_l1035_l1046_l1040_DUPLICATE_6504_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1049_c30_eb5b_return_output;
     -- t8_MUX[uxn_opcodes_h_l1043_c7_f340] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1043_c7_f340_cond <= VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_cond;
     t8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue;
     t8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output := t8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1054_c7_5d8c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1054_c7_5d8c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1046_c7_55cd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1035_c1_8e35] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1054_c7_5d8c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output;

     -- n8_MUX[uxn_opcodes_h_l1046_c7_55cd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1046_c7_55cd_cond <= VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_cond;
     n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue;
     n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output := n8_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1046_c7_55cd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1046_c7_55cd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output := result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1036_c3_dc0e_uxn_opcodes_h_l1036_c3_dc0e_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1035_c1_8e35_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1054_c7_5d8c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;
     -- n8_MUX[uxn_opcodes_h_l1043_c7_f340] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1043_c7_f340_cond <= VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_cond;
     n8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue;
     n8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output := n8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1043_c7_f340] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_return_output := result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;

     -- printf_uxn_opcodes_h_l1036_c3_dc0e[uxn_opcodes_h_l1036_c3_dc0e] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1036_c3_dc0e_uxn_opcodes_h_l1036_c3_dc0e_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1036_c3_dc0e_uxn_opcodes_h_l1036_c3_dc0e_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1043_c7_f340] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1046_c7_55cd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1046_c7_55cd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1043_c7_f340] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1046_c7_55cd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;

     -- t8_MUX[uxn_opcodes_h_l1040_c7_fdab] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond <= VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond;
     t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue;
     t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output := t8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1046_c7_55cd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1040_c7_fdab] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output := result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1040_c7_fdab] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;

     -- t8_MUX[uxn_opcodes_h_l1035_c2_df05] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1035_c2_df05_cond <= VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_cond;
     t8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue;
     t8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output := t8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output;

     -- n8_MUX[uxn_opcodes_h_l1040_c7_fdab] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond <= VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_cond;
     n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue;
     n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output := n8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1040_c7_fdab] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1043_c7_f340] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1043_c7_f340] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1043_c7_f340] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1043_c7_f340_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1035_c2_df05] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_return_output := result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1040_c7_fdab] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1035_c2_df05] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1040_c7_fdab] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1040_c7_fdab] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;

     -- n8_MUX[uxn_opcodes_h_l1035_c2_df05] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1035_c2_df05_cond <= VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_cond;
     n8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue;
     n8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output := n8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1035_c2_df05] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1035_c2_df05_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1040_c7_fdab_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1035_c2_df05] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1035_c2_df05] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1035_c2_df05] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1060_l1031_DUPLICATE_d824 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1060_l1031_DUPLICATE_d824_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8c29(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1035_c2_df05_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1035_c2_df05_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1060_l1031_DUPLICATE_d824_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l1060_l1031_DUPLICATE_d824_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
