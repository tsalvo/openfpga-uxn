-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity inc_0CLK_3045e391 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc_0CLK_3045e391;
architecture arch of inc_0CLK_3045e391 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1437_c6_81c4]
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1437_c1_1825]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1437_c2_5e55]
signal t8_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1437_c2_5e55]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1437_c2_5e55]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1437_c2_5e55]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1437_c2_5e55]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1437_c2_5e55]
signal result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1437_c2_5e55]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l1438_c3_33e3[uxn_opcodes_h_l1438_c3_33e3]
signal printf_uxn_opcodes_h_l1438_c3_33e3_uxn_opcodes_h_l1438_c3_33e3_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1442_c11_d4a1]
signal BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1442_c7_4aed]
signal t8_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1442_c7_4aed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1442_c7_4aed]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1442_c7_4aed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1442_c7_4aed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1442_c7_4aed]
signal result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1442_c7_4aed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1445_c11_15f4]
signal BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1445_c7_3421]
signal t8_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1445_c7_3421]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1445_c7_3421]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1445_c7_3421]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1445_c7_3421]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1445_c7_3421]
signal result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1445_c7_3421]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1448_c32_9555]
signal BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1448_c32_04b2]
signal BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1448_c32_aa09]
signal MUX_uxn_opcodes_h_l1448_c32_aa09_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1448_c32_aa09_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1448_c32_aa09_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1448_c32_aa09_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1450_c11_45a5]
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1450_c7_2ec1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1450_c7_2ec1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1450_c7_2ec1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1450_c7_2ec1]
signal result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1450_c7_2ec1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1454_c24_37a5]
signal BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1456_c11_3268]
signal BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1456_c7_a33f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1456_c7_a33f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_09c5( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.stack_value := ref_toks_5;
      base.is_opc_done := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_left,
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_right,
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_return_output);

-- t8_MUX_uxn_opcodes_h_l1437_c2_5e55
t8_MUX_uxn_opcodes_h_l1437_c2_5e55 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1437_c2_5e55_cond,
t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue,
t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse,
t8_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55
result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55
result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_cond,
result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output);

-- printf_uxn_opcodes_h_l1438_c3_33e3_uxn_opcodes_h_l1438_c3_33e3
printf_uxn_opcodes_h_l1438_c3_33e3_uxn_opcodes_h_l1438_c3_33e3 : entity work.printf_uxn_opcodes_h_l1438_c3_33e3_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1438_c3_33e3_uxn_opcodes_h_l1438_c3_33e3_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1
BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_left,
BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_right,
BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output);

-- t8_MUX_uxn_opcodes_h_l1442_c7_4aed
t8_MUX_uxn_opcodes_h_l1442_c7_4aed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1442_c7_4aed_cond,
t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue,
t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse,
t8_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed
result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed
result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed
result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed
result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_cond,
result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed
result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4
BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_left,
BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_right,
BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output);

-- t8_MUX_uxn_opcodes_h_l1445_c7_3421
t8_MUX_uxn_opcodes_h_l1445_c7_3421 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1445_c7_3421_cond,
t8_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue,
t8_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse,
t8_MUX_uxn_opcodes_h_l1445_c7_3421_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421
result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421
result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421
result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421
result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_cond,
result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421
result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555
BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_left,
BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_right,
BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2
BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_left,
BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_right,
BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_return_output);

-- MUX_uxn_opcodes_h_l1448_c32_aa09
MUX_uxn_opcodes_h_l1448_c32_aa09 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1448_c32_aa09_cond,
MUX_uxn_opcodes_h_l1448_c32_aa09_iftrue,
MUX_uxn_opcodes_h_l1448_c32_aa09_iffalse,
MUX_uxn_opcodes_h_l1448_c32_aa09_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_left,
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_right,
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1
result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1
result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond,
result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5
BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_left,
BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_right,
BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268
BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_left,
BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_right,
BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f
result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f
result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_return_output,
 t8_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output,
 t8_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output,
 t8_MUX_uxn_opcodes_h_l1445_c7_3421_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_return_output,
 MUX_uxn_opcodes_h_l1448_c32_aa09_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1439_c3_22ff : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1438_c3_33e3_uxn_opcodes_h_l1438_c3_33e3_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1443_c3_bf5d : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1453_c3_3518 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_uxn_opcodes_h_l1454_c3_836d : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_1c71_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1450_l1442_l1437_DUPLICATE_48ef_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_eab5_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1450_l1442_l1445_l1437_DUPLICATE_2071_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1450_l1442_l1456_l1445_DUPLICATE_488c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1450_l1445_DUPLICATE_3aae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_09c5_uxn_opcodes_h_l1461_l1433_DUPLICATE_cd6b_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_right := to_unsigned(0, 1);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_right := to_unsigned(128, 8);
     VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1443_c3_bf5d := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1443_c3_bf5d;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1453_c3_3518 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1453_c3_3518;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1439_c3_22ff := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1439_c3_22ff;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_right := to_unsigned(3, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1450_c11_45a5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l1448_c32_9555] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_left;
     BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_return_output := BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1450_l1445_DUPLICATE_3aae LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1450_l1445_DUPLICATE_3aae_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1450_l1442_l1437_DUPLICATE_48ef LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1450_l1442_l1437_DUPLICATE_48ef_return_output := result.is_sp_shift;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_eab5 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_eab5_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1442_c11_d4a1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_1c71 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_1c71_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1437_c6_81c4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1445_c11_15f4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1456_c11_3268] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_left;
     BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_return_output := BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1454_c24_37a5] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1450_l1442_l1445_l1437_DUPLICATE_2071 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1450_l1442_l1445_l1437_DUPLICATE_2071_return_output := result.stack_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1450_l1442_l1456_l1445_DUPLICATE_488c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1450_l1442_l1456_l1445_DUPLICATE_488c_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1448_c32_9555_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_81c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1442_c11_d4a1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1445_c11_15f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_45a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1456_c11_3268_return_output;
     VAR_result_stack_value_uxn_opcodes_h_l1454_c3_836d := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1454_c24_37a5_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_eab5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_eab5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1442_l1445_l1437_DUPLICATE_eab5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1450_l1442_l1456_l1445_DUPLICATE_488c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1450_l1442_l1456_l1445_DUPLICATE_488c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1450_l1442_l1456_l1445_DUPLICATE_488c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1450_l1442_l1456_l1445_DUPLICATE_488c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1450_l1442_l1437_DUPLICATE_48ef_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1450_l1442_l1437_DUPLICATE_48ef_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1450_l1442_l1437_DUPLICATE_48ef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_1c71_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_1c71_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_1c71_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1442_l1456_l1445_l1437_DUPLICATE_1c71_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1450_l1445_DUPLICATE_3aae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1450_l1445_DUPLICATE_3aae_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1450_l1442_l1445_l1437_DUPLICATE_2071_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1450_l1442_l1445_l1437_DUPLICATE_2071_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1450_l1442_l1445_l1437_DUPLICATE_2071_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1450_l1442_l1445_l1437_DUPLICATE_2071_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue := VAR_result_stack_value_uxn_opcodes_h_l1454_c3_836d;
     -- result_stack_value_MUX[uxn_opcodes_h_l1450_c7_2ec1] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output := result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1456_c7_a33f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1437_c1_1825] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1450_c7_2ec1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1448_c32_04b2] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_left;
     BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_return_output := BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1456_c7_a33f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1445_c7_3421] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1445_c7_3421_cond <= VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_cond;
     t8_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue;
     t8_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_return_output := t8_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1450_c7_2ec1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1448_c32_04b2_return_output;
     VAR_printf_uxn_opcodes_h_l1438_c3_33e3_uxn_opcodes_h_l1438_c3_33e3_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1437_c1_1825_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1456_c7_a33f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l1445_c7_3421] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_return_output := result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1450_c7_2ec1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1450_c7_2ec1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output;

     -- t8_MUX[uxn_opcodes_h_l1442_c7_4aed] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1442_c7_4aed_cond <= VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_cond;
     t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue;
     t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output := t8_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1445_c7_3421] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;

     -- MUX[uxn_opcodes_h_l1448_c32_aa09] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1448_c32_aa09_cond <= VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_cond;
     MUX_uxn_opcodes_h_l1448_c32_aa09_iftrue <= VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_iftrue;
     MUX_uxn_opcodes_h_l1448_c32_aa09_iffalse <= VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_return_output := MUX_uxn_opcodes_h_l1448_c32_aa09_return_output;

     -- printf_uxn_opcodes_h_l1438_c3_33e3[uxn_opcodes_h_l1438_c3_33e3] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1438_c3_33e3_uxn_opcodes_h_l1438_c3_33e3_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1438_c3_33e3_uxn_opcodes_h_l1438_c3_33e3_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1445_c7_3421] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue := VAR_MUX_uxn_opcodes_h_l1448_c32_aa09_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_2ec1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;
     -- t8_MUX[uxn_opcodes_h_l1437_c2_5e55] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1437_c2_5e55_cond <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_cond;
     t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue;
     t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output := t8_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1442_c7_4aed] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output := result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1445_c7_3421] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1445_c7_3421] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1445_c7_3421] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1442_c7_4aed] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1442_c7_4aed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1445_c7_3421_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l1437_c2_5e55] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output := result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1442_c7_4aed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1437_c2_5e55] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1442_c7_4aed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1442_c7_4aed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1437_c2_5e55] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1442_c7_4aed_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1437_c2_5e55] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1437_c2_5e55] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1437_c2_5e55] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_09c5_uxn_opcodes_h_l1461_l1433_DUPLICATE_cd6b LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_09c5_uxn_opcodes_h_l1461_l1433_DUPLICATE_cd6b_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_09c5(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_5e55_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_09c5_uxn_opcodes_h_l1461_l1433_DUPLICATE_cd6b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_09c5_uxn_opcodes_h_l1461_l1433_DUPLICATE_cd6b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
