-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity add_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end add_0CLK_fedec265;
architecture arch of add_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l857_c6_864a]
signal BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l857_c2_5dc0]
signal n8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l857_c2_5dc0]
signal t8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l857_c2_5dc0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l857_c2_5dc0]
signal result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l857_c2_5dc0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l857_c2_5dc0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l857_c2_5dc0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l857_c2_5dc0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l862_c11_2af8]
signal BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l862_c7_92f2]
signal n8_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l862_c7_92f2]
signal t8_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l862_c7_92f2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l862_c7_92f2]
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l862_c7_92f2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l862_c7_92f2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l862_c7_92f2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l862_c7_92f2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l865_c11_d9cf]
signal BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l865_c7_5833]
signal n8_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l865_c7_5833]
signal t8_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l865_c7_5833]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l865_c7_5833]
signal result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l865_c7_5833]
signal result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l865_c7_5833]
signal result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l865_c7_5833]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l865_c7_5833]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l869_c11_a113]
signal BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l869_c7_1e7e]
signal n8_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l869_c7_1e7e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l869_c7_1e7e]
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l869_c7_1e7e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l869_c7_1e7e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l869_c7_1e7e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l869_c7_1e7e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l872_c11_b097]
signal BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l872_c7_29ce]
signal n8_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l872_c7_29ce]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l872_c7_29ce]
signal result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l872_c7_29ce]
signal result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l872_c7_29ce]
signal result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l872_c7_29ce]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l872_c7_29ce]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l875_c30_feef]
signal sp_relative_shift_uxn_opcodes_h_l875_c30_feef_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l875_c30_feef_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l875_c30_feef_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l875_c30_feef_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l878_c21_c322]
signal BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_right : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l880_c11_b232]
signal BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l880_c7_6ce5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l880_c7_6ce5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l880_c7_6ce5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a
BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_left,
BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_right,
BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output);

-- n8_MUX_uxn_opcodes_h_l857_c2_5dc0
n8_MUX_uxn_opcodes_h_l857_c2_5dc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond,
n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue,
n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse,
n8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output);

-- t8_MUX_uxn_opcodes_h_l857_c2_5dc0
t8_MUX_uxn_opcodes_h_l857_c2_5dc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond,
t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue,
t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse,
t8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0
result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_cond,
result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0
result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0
result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0
result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0
result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8
BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_left,
BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_right,
BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output);

-- n8_MUX_uxn_opcodes_h_l862_c7_92f2
n8_MUX_uxn_opcodes_h_l862_c7_92f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l862_c7_92f2_cond,
n8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue,
n8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse,
n8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output);

-- t8_MUX_uxn_opcodes_h_l862_c7_92f2
t8_MUX_uxn_opcodes_h_l862_c7_92f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l862_c7_92f2_cond,
t8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue,
t8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse,
t8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2
result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_cond,
result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf
BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_left,
BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_right,
BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output);

-- n8_MUX_uxn_opcodes_h_l865_c7_5833
n8_MUX_uxn_opcodes_h_l865_c7_5833 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l865_c7_5833_cond,
n8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue,
n8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse,
n8_MUX_uxn_opcodes_h_l865_c7_5833_return_output);

-- t8_MUX_uxn_opcodes_h_l865_c7_5833
t8_MUX_uxn_opcodes_h_l865_c7_5833 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l865_c7_5833_cond,
t8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue,
t8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse,
t8_MUX_uxn_opcodes_h_l865_c7_5833_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833
result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_cond,
result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833
result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833
result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833
result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833
result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113
BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_left,
BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_right,
BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output);

-- n8_MUX_uxn_opcodes_h_l869_c7_1e7e
n8_MUX_uxn_opcodes_h_l869_c7_1e7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l869_c7_1e7e_cond,
n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue,
n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse,
n8_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e
result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_cond,
result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097
BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_left,
BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_right,
BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output);

-- n8_MUX_uxn_opcodes_h_l872_c7_29ce
n8_MUX_uxn_opcodes_h_l872_c7_29ce : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l872_c7_29ce_cond,
n8_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue,
n8_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse,
n8_MUX_uxn_opcodes_h_l872_c7_29ce_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce
result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_cond,
result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce
result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce
result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce
result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce
result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output);

-- sp_relative_shift_uxn_opcodes_h_l875_c30_feef
sp_relative_shift_uxn_opcodes_h_l875_c30_feef : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l875_c30_feef_ins,
sp_relative_shift_uxn_opcodes_h_l875_c30_feef_x,
sp_relative_shift_uxn_opcodes_h_l875_c30_feef_y,
sp_relative_shift_uxn_opcodes_h_l875_c30_feef_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322
BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322 : entity work.BIN_OP_PLUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_left,
BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_right,
BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232
BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_left,
BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_right,
BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5
result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5
result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5
result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output,
 n8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
 t8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output,
 n8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output,
 t8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output,
 n8_MUX_uxn_opcodes_h_l865_c7_5833_return_output,
 t8_MUX_uxn_opcodes_h_l865_c7_5833_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output,
 n8_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output,
 n8_MUX_uxn_opcodes_h_l872_c7_29ce_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output,
 sp_relative_shift_uxn_opcodes_h_l875_c30_feef_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l859_c3_f7d0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l863_c3_e009 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l867_c3_5a9e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l870_c3_2bd1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l877_c3_291f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l872_c7_29ce_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l878_c3_d70b : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_558a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_765b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_35a3_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_7c51_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l869_l865_l862_l880_l872_DUPLICATE_bd7d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l886_l853_DUPLICATE_2b03_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l867_c3_5a9e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l867_c3_5a9e;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l859_c3_f7d0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l859_c3_f7d0;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l877_c3_291f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l877_c3_291f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l863_c3_e009 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l863_c3_e009;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l870_c3_2bd1 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l870_c3_2bd1;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l869_c11_a113] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_left;
     BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output := BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l872_c11_b097] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_left;
     BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output := BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l865_c11_d9cf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_left;
     BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output := BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l872_c7_29ce] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l872_c7_29ce_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_765b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_765b_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l862_c11_2af8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_left;
     BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output := BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l869_l865_l862_l880_l872_DUPLICATE_bd7d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l869_l865_l862_l880_l872_DUPLICATE_bd7d_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l857_c6_864a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_left;
     BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output := BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l880_c11_b232] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_left;
     BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_return_output := BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_558a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_558a_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_7c51 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_7c51_return_output := result.is_sp_shift;

     -- BIN_OP_PLUS[uxn_opcodes_h_l878_c21_c322] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_left;
     BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_return_output := BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_35a3 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_35a3_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l875_c30_feef] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l875_c30_feef_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_ins;
     sp_relative_shift_uxn_opcodes_h_l875_c30_feef_x <= VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_x;
     sp_relative_shift_uxn_opcodes_h_l875_c30_feef_y <= VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_return_output := sp_relative_shift_uxn_opcodes_h_l875_c30_feef_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l857_c6_864a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_2af8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l865_c11_d9cf_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_a113_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l872_c11_b097_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l880_c11_b232_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l878_c3_d70b := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l878_c21_c322_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_35a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_35a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_35a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_35a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_35a3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l869_l865_l862_l880_l872_DUPLICATE_bd7d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l869_l865_l862_l880_l872_DUPLICATE_bd7d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l869_l865_l862_l880_l872_DUPLICATE_bd7d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l869_l865_l862_l880_l872_DUPLICATE_bd7d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l869_l865_l862_l880_l872_DUPLICATE_bd7d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_7c51_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_7c51_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_7c51_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_7c51_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_7c51_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_765b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_765b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_765b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_765b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l869_l865_l862_l857_l880_DUPLICATE_765b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_558a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_558a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_558a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_558a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l869_l865_l862_l857_l872_DUPLICATE_558a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l872_c7_29ce_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l875_c30_feef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue := VAR_result_u8_value_uxn_opcodes_h_l878_c3_d70b;
     -- n8_MUX[uxn_opcodes_h_l872_c7_29ce] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l872_c7_29ce_cond <= VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_cond;
     n8_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue;
     n8_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_return_output := n8_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;

     -- t8_MUX[uxn_opcodes_h_l865_c7_5833] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l865_c7_5833_cond <= VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_cond;
     t8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue;
     t8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_return_output := t8_MUX_uxn_opcodes_h_l865_c7_5833_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l880_c7_6ce5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l872_c7_29ce] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l872_c7_29ce] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l880_c7_6ce5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l872_c7_29ce] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_cond;
     result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_return_output := result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l880_c7_6ce5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l880_c7_6ce5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l865_c7_5833_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l872_c7_29ce] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l872_c7_29ce] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;

     -- n8_MUX[uxn_opcodes_h_l869_c7_1e7e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l869_c7_1e7e_cond <= VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_cond;
     n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue;
     n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output := n8_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l869_c7_1e7e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l872_c7_29ce] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;

     -- t8_MUX[uxn_opcodes_h_l862_c7_92f2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l862_c7_92f2_cond <= VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_cond;
     t8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue;
     t8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output := t8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l869_c7_1e7e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output := result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l869_c7_1e7e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse := VAR_n8_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l872_c7_29ce_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l869_c7_1e7e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;

     -- n8_MUX[uxn_opcodes_h_l865_c7_5833] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l865_c7_5833_cond <= VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_cond;
     n8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_iftrue;
     n8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_return_output := n8_MUX_uxn_opcodes_h_l865_c7_5833_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l865_c7_5833] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l869_c7_1e7e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l865_c7_5833] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_cond;
     result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_return_output := result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_return_output;

     -- t8_MUX[uxn_opcodes_h_l857_c2_5dc0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond <= VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond;
     t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue;
     t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output := t8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l865_c7_5833] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l869_c7_1e7e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l865_c7_5833_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_1e7e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l865_c7_5833_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l865_c7_5833_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l865_c7_5833] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l865_c7_5833] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l862_c7_92f2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_return_output := result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l862_c7_92f2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l865_c7_5833] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_return_output;

     -- n8_MUX[uxn_opcodes_h_l862_c7_92f2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l862_c7_92f2_cond <= VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_cond;
     n8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue;
     n8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output := n8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l862_c7_92f2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l865_c7_5833_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l865_c7_5833_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l865_c7_5833_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l862_c7_92f2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l857_c2_5dc0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output;

     -- n8_MUX[uxn_opcodes_h_l857_c2_5dc0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond <= VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_cond;
     n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue;
     n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output := n8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l857_c2_5dc0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l862_c7_92f2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l857_c2_5dc0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output := result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l862_c7_92f2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_92f2_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l857_c2_5dc0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l857_c2_5dc0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l857_c2_5dc0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l886_l853_DUPLICATE_2b03 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l886_l853_DUPLICATE_2b03_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l857_c2_5dc0_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l886_l853_DUPLICATE_2b03_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l886_l853_DUPLICATE_2b03_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
