-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity sth_0CLK_edc09f97 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_edc09f97;
architecture arch of sth_0CLK_edc09f97 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2777_c6_6865]
signal BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2777_c1_c50f]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2777_c2_a0a6]
signal t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2777_c2_a0a6]
signal result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2777_c2_a0a6]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2777_c2_a0a6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2777_c2_a0a6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : signed(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2777_c2_a0a6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2777_c2_a0a6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2777_c2_a0a6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2777_c2_a0a6]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l2778_c3_a53f[uxn_opcodes_h_l2778_c3_a53f]
signal printf_uxn_opcodes_h_l2778_c3_a53f_uxn_opcodes_h_l2778_c3_a53f_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2783_c11_0109]
signal BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2783_c7_c8c8]
signal t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2783_c7_c8c8]
signal result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2783_c7_c8c8]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2783_c7_c8c8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2783_c7_c8c8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : signed(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2783_c7_c8c8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2783_c7_c8c8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2783_c7_c8c8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2783_c7_c8c8]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2786_c11_0e33]
signal BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2786_c7_b231]
signal t8_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2786_c7_b231]
signal result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2786_c7_b231]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2786_c7_b231]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2786_c7_b231]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : signed(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2786_c7_b231]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2786_c7_b231]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2786_c7_b231]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(0 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2786_c7_b231]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2790_c32_889f]
signal BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l2790_c32_7f59]
signal BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2790_c32_d122]
signal MUX_uxn_opcodes_h_l2790_c32_d122_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2790_c32_d122_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2790_c32_d122_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2790_c32_d122_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2792_c11_91b4]
signal BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2792_c7_bde6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2792_c7_bde6]
signal result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2792_c7_bde6]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2792_c7_bde6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2792_c7_bde6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : signed(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2792_c7_bde6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2792_c7_bde6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2796_c11_281c]
signal BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2796_c7_3e2a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2796_c7_3e2a]
signal result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2796_c7_3e2a]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2796_c7_3e2a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2796_c7_3e2a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2796_c7_3e2a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2802_c11_211e]
signal BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2802_c7_df5d]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2802_c7_df5d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2802_c7_df5d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c029( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_value := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_sp_shift := ref_toks_6;
      base.is_opc_done := ref_toks_7;
      base.is_stack_read := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865
BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_left,
BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_right,
BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_return_output);

-- t8_MUX_uxn_opcodes_h_l2777_c2_a0a6
t8_MUX_uxn_opcodes_h_l2777_c2_a0a6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond,
t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue,
t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse,
t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6
result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond,
result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6
result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6
result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6
result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6
result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output);

-- printf_uxn_opcodes_h_l2778_c3_a53f_uxn_opcodes_h_l2778_c3_a53f
printf_uxn_opcodes_h_l2778_c3_a53f_uxn_opcodes_h_l2778_c3_a53f : entity work.printf_uxn_opcodes_h_l2778_c3_a53f_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2778_c3_a53f_uxn_opcodes_h_l2778_c3_a53f_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109
BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_left,
BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_right,
BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output);

-- t8_MUX_uxn_opcodes_h_l2783_c7_c8c8
t8_MUX_uxn_opcodes_h_l2783_c7_c8c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond,
t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue,
t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse,
t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8
result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond,
result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8
result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8
result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8
result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8
result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33
BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_left,
BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_right,
BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output);

-- t8_MUX_uxn_opcodes_h_l2786_c7_b231
t8_MUX_uxn_opcodes_h_l2786_c7_b231 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2786_c7_b231_cond,
t8_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue,
t8_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse,
t8_MUX_uxn_opcodes_h_l2786_c7_b231_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231
result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_cond,
result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231
result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231
result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231
result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231
result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231
result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f
BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_left,
BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_right,
BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59
BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_left,
BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_right,
BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_return_output);

-- MUX_uxn_opcodes_h_l2790_c32_d122
MUX_uxn_opcodes_h_l2790_c32_d122 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2790_c32_d122_cond,
MUX_uxn_opcodes_h_l2790_c32_d122_iftrue,
MUX_uxn_opcodes_h_l2790_c32_d122_iffalse,
MUX_uxn_opcodes_h_l2790_c32_d122_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4
BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_left,
BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_right,
BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6
result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6
result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_cond,
result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6
result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6
result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c
BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_left,
BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_right,
BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a
result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a
result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond,
result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a
result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a
result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e
BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_left,
BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_right,
BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d
result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d
result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_return_output,
 t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output,
 t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output,
 t8_MUX_uxn_opcodes_h_l2786_c7_b231_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_return_output,
 BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_return_output,
 MUX_uxn_opcodes_h_l2790_c32_d122_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2780_c3_0e53 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2778_c3_a53f_uxn_opcodes_h_l2778_c3_a53f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2784_c3_f77c : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2790_c32_d122_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2790_c32_d122_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2790_c32_d122_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2790_c32_d122_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2794_c3_8b47 : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2799_c3_7941 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2796_l2792_l2786_l2783_l2777_DUPLICATE_92c8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2802_l2796_l2786_l2783_l2777_DUPLICATE_ee5b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2802_l2792_l2786_l2783_l2777_DUPLICATE_aa8e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2783_l2777_l2792_DUPLICATE_85d0_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2783_l2796_l2777_l2792_DUPLICATE_c378_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2802_l2796_l2792_l2786_l2783_DUPLICATE_ab5a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2783_l2786_DUPLICATE_cac1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2796_l2786_l2792_DUPLICATE_1dfb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c029_uxn_opcodes_h_l2773_l2808_DUPLICATE_e05e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l2790_c32_d122_iffalse := resize(to_signed(-1, 2), 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2780_c3_0e53 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2780_c3_0e53;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_right := to_unsigned(5, 3);
     VAR_MUX_uxn_opcodes_h_l2790_c32_d122_iftrue := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2794_c3_8b47 := signed(std_logic_vector(resize(to_unsigned(2, 2), 8)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2794_c3_8b47;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_right := to_unsigned(3, 2);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2799_c3_7941 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2799_c3_7941;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2784_c3_f77c := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2784_c3_f77c;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_right := to_unsigned(128, 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2796_l2786_l2792_DUPLICATE_1dfb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2796_l2786_l2792_DUPLICATE_1dfb_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2783_l2777_l2792_DUPLICATE_85d0 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2783_l2777_l2792_DUPLICATE_85d0_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2802_c11_211e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2783_l2796_l2777_l2792_DUPLICATE_c378 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2783_l2796_l2777_l2792_DUPLICATE_c378_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2802_l2796_l2786_l2783_l2777_DUPLICATE_ee5b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2802_l2796_l2786_l2783_l2777_DUPLICATE_ee5b_return_output := result.is_stack_index_flipped;

     -- BIN_OP_AND[uxn_opcodes_h_l2790_c32_889f] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_left;
     BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_return_output := BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2802_l2792_l2786_l2783_l2777_DUPLICATE_aa8e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2802_l2792_l2786_l2783_l2777_DUPLICATE_aa8e_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2802_l2796_l2792_l2786_l2783_DUPLICATE_ab5a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2802_l2796_l2792_l2786_l2783_DUPLICATE_ab5a_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2786_c11_0e33] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_left;
     BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output := BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2792_c11_91b4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2783_l2786_DUPLICATE_cac1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2783_l2786_DUPLICATE_cac1_return_output := result.is_stack_read;

     -- BIN_OP_EQ[uxn_opcodes_h_l2777_c6_6865] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_left;
     BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output := BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2783_c11_0109] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_left;
     BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output := BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2796_c11_281c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2796_l2792_l2786_l2783_l2777_DUPLICATE_92c8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2796_l2792_l2786_l2783_l2777_DUPLICATE_92c8_return_output := result.stack_value;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_left := VAR_BIN_OP_AND_uxn_opcodes_h_l2790_c32_889f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2777_c6_6865_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2783_c11_0109_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2786_c11_0e33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2792_c11_91b4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2796_c11_281c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2802_c11_211e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2783_l2777_l2792_DUPLICATE_85d0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2783_l2777_l2792_DUPLICATE_85d0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2783_l2777_l2792_DUPLICATE_85d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2802_l2796_l2792_l2786_l2783_DUPLICATE_ab5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2802_l2796_l2792_l2786_l2783_DUPLICATE_ab5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2802_l2796_l2792_l2786_l2783_DUPLICATE_ab5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2802_l2796_l2792_l2786_l2783_DUPLICATE_ab5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2802_l2796_l2792_l2786_l2783_DUPLICATE_ab5a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2783_l2796_l2777_l2792_DUPLICATE_c378_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2783_l2796_l2777_l2792_DUPLICATE_c378_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2783_l2796_l2777_l2792_DUPLICATE_c378_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2783_l2796_l2777_l2792_DUPLICATE_c378_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2802_l2796_l2786_l2783_l2777_DUPLICATE_ee5b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2802_l2796_l2786_l2783_l2777_DUPLICATE_ee5b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2802_l2796_l2786_l2783_l2777_DUPLICATE_ee5b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2802_l2796_l2786_l2783_l2777_DUPLICATE_ee5b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2802_l2796_l2786_l2783_l2777_DUPLICATE_ee5b_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2783_l2786_DUPLICATE_cac1_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2783_l2786_DUPLICATE_cac1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2802_l2792_l2786_l2783_l2777_DUPLICATE_aa8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2802_l2792_l2786_l2783_l2777_DUPLICATE_aa8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2802_l2792_l2786_l2783_l2777_DUPLICATE_aa8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2802_l2792_l2786_l2783_l2777_DUPLICATE_aa8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2802_l2792_l2786_l2783_l2777_DUPLICATE_aa8e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2796_l2786_l2792_DUPLICATE_1dfb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2796_l2786_l2792_DUPLICATE_1dfb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2796_l2786_l2792_DUPLICATE_1dfb_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2796_l2792_l2786_l2783_l2777_DUPLICATE_92c8_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2796_l2792_l2786_l2783_l2777_DUPLICATE_92c8_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2796_l2792_l2786_l2783_l2777_DUPLICATE_92c8_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2796_l2792_l2786_l2783_l2777_DUPLICATE_92c8_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2796_l2792_l2786_l2783_l2777_DUPLICATE_92c8_return_output;
     -- BIN_OP_GT[uxn_opcodes_h_l2790_c32_7f59] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_left;
     BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_return_output := BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2802_c7_df5d] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2802_c7_df5d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2802_c7_df5d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output;

     -- t8_MUX[uxn_opcodes_h_l2786_c7_b231] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2786_c7_b231_cond <= VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_cond;
     t8_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue;
     t8_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_return_output := t8_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2796_c7_3e2a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2796_c7_3e2a] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output := result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2796_c7_3e2a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2786_c7_b231] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2792_c7_bde6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2777_c1_c50f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l2790_c32_d122_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l2790_c32_7f59_return_output;
     VAR_printf_uxn_opcodes_h_l2778_c3_a53f_uxn_opcodes_h_l2778_c3_a53f_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2777_c1_c50f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2802_c7_df5d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2792_c7_bde6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2796_c7_3e2a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2792_c7_bde6] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output := result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;

     -- t8_MUX[uxn_opcodes_h_l2783_c7_c8c8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond <= VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond;
     t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue;
     t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output := t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2783_c7_c8c8] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;

     -- MUX[uxn_opcodes_h_l2790_c32_d122] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2790_c32_d122_cond <= VAR_MUX_uxn_opcodes_h_l2790_c32_d122_cond;
     MUX_uxn_opcodes_h_l2790_c32_d122_iftrue <= VAR_MUX_uxn_opcodes_h_l2790_c32_d122_iftrue;
     MUX_uxn_opcodes_h_l2790_c32_d122_iffalse <= VAR_MUX_uxn_opcodes_h_l2790_c32_d122_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2790_c32_d122_return_output := MUX_uxn_opcodes_h_l2790_c32_d122_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2796_c7_3e2a] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;

     -- printf_uxn_opcodes_h_l2778_c3_a53f[uxn_opcodes_h_l2778_c3_a53f] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2778_c3_a53f_uxn_opcodes_h_l2778_c3_a53f_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2778_c3_a53f_uxn_opcodes_h_l2778_c3_a53f_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2796_c7_3e2a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2792_c7_bde6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue := VAR_MUX_uxn_opcodes_h_l2790_c32_d122_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2796_c7_3e2a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2792_c7_bde6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;

     -- t8_MUX[uxn_opcodes_h_l2777_c2_a0a6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond <= VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond;
     t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue;
     t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output := t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2786_c7_b231] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_return_output := result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2786_c7_b231] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2786_c7_b231] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2786_c7_b231] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2792_c7_bde6] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2792_c7_bde6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2777_c2_a0a6] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2792_c7_bde6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output;
     -- result_stack_value_MUX[uxn_opcodes_h_l2783_c7_c8c8] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output := result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2783_c7_c8c8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2786_c7_b231] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2786_c7_b231] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2786_c7_b231] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2783_c7_c8c8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2783_c7_c8c8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2786_c7_b231_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2783_c7_c8c8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2777_c2_a0a6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2783_c7_c8c8] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2783_c7_c8c8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2777_c2_a0a6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2777_c2_a0a6] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output := result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2777_c2_a0a6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2783_c7_c8c8_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2777_c2_a0a6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2777_c2_a0a6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2777_c2_a0a6] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c029_uxn_opcodes_h_l2773_l2808_DUPLICATE_e05e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c029_uxn_opcodes_h_l2773_l2808_DUPLICATE_e05e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c029(
     result,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2777_c2_a0a6_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c029_uxn_opcodes_h_l2773_l2808_DUPLICATE_e05e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c029_uxn_opcodes_h_l2773_l2808_DUPLICATE_e05e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
