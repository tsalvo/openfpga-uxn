-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 42
entity jci_0CLK_4351dde2 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jci_0CLK_4351dde2;
architecture arch of jci_0CLK_4351dde2 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l71_c6_3881]
signal BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l71_c2_beb1]
signal tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(15 downto 0);

-- t8_MUX[uxn_opcodes_h_l71_c2_beb1]
signal t8_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l71_c2_beb1]
signal result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l71_c2_beb1]
signal result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l71_c2_beb1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l71_c2_beb1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l71_c2_beb1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l71_c2_beb1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l71_c2_beb1]
signal result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l71_c2_beb1]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l71_c2_beb1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l85_c11_d121]
signal BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l85_c7_2701]
signal tmp16_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(15 downto 0);

-- t8_MUX[uxn_opcodes_h_l85_c7_2701]
signal t8_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l85_c7_2701]
signal result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l85_c7_2701]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l85_c7_2701]
signal result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l85_c7_2701]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l85_c7_2701]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l88_c22_e57e]
signal BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l90_c11_4e7b]
signal BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l90_c7_7d27]
signal tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : unsigned(15 downto 0);

-- t8_MUX[uxn_opcodes_h_l90_c7_7d27]
signal t8_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l90_c7_7d27]
signal result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l90_c7_7d27]
signal result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l90_c7_7d27]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l90_c7_7d27]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : signed(3 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l93_c3_cfb0]
signal CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l96_c11_c4ea]
signal BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l96_c7_2fa9]
signal tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l96_c7_2fa9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l96_c7_2fa9]
signal result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l96_c7_2fa9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output : unsigned(0 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l97_c3_1523]
signal BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l99_c22_cfef]
signal BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l99_c32_792b]
signal BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_right : unsigned(1 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_return_output : unsigned(16 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l99_c42_fe5d]
signal BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_right : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_return_output : unsigned(16 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l99_c42_bc76]
signal BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_left : unsigned(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_right : unsigned(1 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_return_output : unsigned(17 downto 0);

-- MUX[uxn_opcodes_h_l99_c22_e9ee]
signal MUX_uxn_opcodes_h_l99_c22_e9ee_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l99_c22_e9ee_iftrue : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l99_c22_e9ee_iffalse : unsigned(15 downto 0);
signal MUX_uxn_opcodes_h_l99_c22_e9ee_return_output : unsigned(15 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_161f( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_vram_write := ref_toks_1;
      base.u16_value := ref_toks_2;
      base.is_pc_updated := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.sp_relative_shift := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881
BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_left,
BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_right,
BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output);

-- tmp16_MUX_uxn_opcodes_h_l71_c2_beb1
tmp16_MUX_uxn_opcodes_h_l71_c2_beb1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_cond,
tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue,
tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse,
tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

-- t8_MUX_uxn_opcodes_h_l71_c2_beb1
t8_MUX_uxn_opcodes_h_l71_c2_beb1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l71_c2_beb1_cond,
t8_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue,
t8_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse,
t8_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1
result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1
result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_cond,
result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1
result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1
result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1
result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1
result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1
result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121
BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_left,
BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_right,
BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output);

-- tmp16_MUX_uxn_opcodes_h_l85_c7_2701
tmp16_MUX_uxn_opcodes_h_l85_c7_2701 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l85_c7_2701_cond,
tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iftrue,
tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iffalse,
tmp16_MUX_uxn_opcodes_h_l85_c7_2701_return_output);

-- t8_MUX_uxn_opcodes_h_l85_c7_2701
t8_MUX_uxn_opcodes_h_l85_c7_2701 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l85_c7_2701_cond,
t8_MUX_uxn_opcodes_h_l85_c7_2701_iftrue,
t8_MUX_uxn_opcodes_h_l85_c7_2701_iffalse,
t8_MUX_uxn_opcodes_h_l85_c7_2701_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701
result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_cond,
result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701
result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701
result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701
result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e
BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_left,
BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_right,
BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b
BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_left,
BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_right,
BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output);

-- tmp16_MUX_uxn_opcodes_h_l90_c7_7d27
tmp16_MUX_uxn_opcodes_h_l90_c7_7d27 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_cond,
tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue,
tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse,
tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_return_output);

-- t8_MUX_uxn_opcodes_h_l90_c7_7d27
t8_MUX_uxn_opcodes_h_l90_c7_7d27 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l90_c7_7d27_cond,
t8_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue,
t8_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse,
t8_MUX_uxn_opcodes_h_l90_c7_7d27_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27
result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27
result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_cond,
result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27
result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27
result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_return_output);

-- CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0
CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_x,
CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea
BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_left,
BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_right,
BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_return_output);

-- tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9
tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_cond,
tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue,
tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse,
tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9
result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9
result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_cond,
result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9
result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l97_c3_1523
BIN_OP_OR_uxn_opcodes_h_l97_c3_1523 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_left,
BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_right,
BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef
BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_left,
BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_right,
BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b
BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b : entity work.BIN_OP_PLUS_uint16_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_left,
BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_right,
BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d
BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d : entity work.BIN_OP_PLUS_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_left,
BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_right,
BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76
BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76 : entity work.BIN_OP_PLUS_uint17_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_left,
BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_right,
BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_return_output);

-- MUX_uxn_opcodes_h_l99_c22_e9ee
MUX_uxn_opcodes_h_l99_c22_e9ee : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l99_c22_e9ee_cond,
MUX_uxn_opcodes_h_l99_c22_e9ee_iftrue,
MUX_uxn_opcodes_h_l99_c22_e9ee_iffalse,
MUX_uxn_opcodes_h_l99_c22_e9ee_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 tmp16,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output,
 tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
 t8_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output,
 tmp16_MUX_uxn_opcodes_h_l85_c7_2701_return_output,
 t8_MUX_uxn_opcodes_h_l85_c7_2701_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output,
 tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_return_output,
 t8_MUX_uxn_opcodes_h_l90_c7_7d27_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_return_output,
 CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_return_output,
 tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output,
 BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_return_output,
 MUX_uxn_opcodes_h_l99_c22_e9ee_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l81_c3_fede : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l76_c3_ac45 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l88_c3_b381 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l86_c3_64ad : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l85_c7_2701_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l87_c3_83f2 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l94_c3_4bf5 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l90_c7_7d27_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_return_output : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_iftrue : unsigned(15 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_iffalse : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_left : unsigned(16 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_return_output : unsigned(17 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_6e0f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_618e_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l92_l97_DUPLICATE_2d2c_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l90_l96_DUPLICATE_7057_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_161f_uxn_opcodes_h_l103_l66_DUPLICATE_39ef_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp16 := tmp16;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l76_c3_ac45 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l76_c3_ac45;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l94_c3_4bf5 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l94_c3_4bf5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l87_c3_83f2 := resize(to_signed(-1, 2), 4);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l87_c3_83f2;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l81_c3_fede := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l81_c3_fede;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_right := to_unsigned(2, 2);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l86_c3_64ad := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l86_c3_64ad;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_left := VAR_pc;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_left := VAR_pc;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_left := VAR_pc;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse := t8;
     VAR_BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_left := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse := tmp16;
     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l90_c7_7d27] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l90_c7_7d27_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l96_c11_c4ea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_left;
     BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_return_output := BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l99_c22_cfef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_left;
     BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_return_output := BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_618e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_618e_return_output := result.is_opc_done;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l92_l97_DUPLICATE_2d2c LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l92_l97_DUPLICATE_2d2c_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_ram_read);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_6e0f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_6e0f_return_output := result.is_pc_updated;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l71_c2_beb1_return_output := result.is_vram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l71_c2_beb1_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l90_c11_4e7b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_left;
     BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output := BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l71_c2_beb1_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l85_c11_d121] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_left;
     BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output := BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l71_c6_3881] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_left;
     BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output := BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l85_c7_2701] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l85_c7_2701_return_output := result.stack_address_sp_offset;

     -- BIN_OP_PLUS[uxn_opcodes_h_l88_c22_e57e] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_left;
     BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_return_output := BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l90_l96_DUPLICATE_7057 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l90_l96_DUPLICATE_7057_return_output := result.u16_value;

     -- BIN_OP_PLUS[uxn_opcodes_h_l99_c32_792b] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_left;
     BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_return_output := BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_return_output;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l71_c2_beb1_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l71_c6_3881_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l85_c11_d121_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l90_c11_4e7b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l96_c11_c4ea_return_output;
     VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l99_c22_cfef_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l88_c3_b381 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l88_c22_e57e_return_output, 16);
     VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_iftrue := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c32_792b_return_output, 16);
     VAR_BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l92_l97_DUPLICATE_2d2c_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l92_l97_DUPLICATE_2d2c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l90_l96_DUPLICATE_7057_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l90_l96_DUPLICATE_7057_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_618e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_618e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_618e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_6e0f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_6e0f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l90_l96_l85_DUPLICATE_6e0f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l71_c2_beb1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l71_c2_beb1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l71_c2_beb1_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l71_c2_beb1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l90_c7_7d27_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l85_c7_2701_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iftrue := VAR_result_u16_value_uxn_opcodes_h_l88_c3_b381;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l90_c7_7d27] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l97_c3_1523] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_left;
     BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_return_output := BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l96_c7_2fa9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output;

     -- t8_MUX[uxn_opcodes_h_l90_c7_7d27] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l90_c7_7d27_cond <= VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_cond;
     t8_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue;
     t8_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_return_output := t8_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l96_c7_2fa9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l85_c7_2701] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l93_c3_cfb0] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_x <= VAR_CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_return_output := CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;

     -- Submodule level 2
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_right := VAR_BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l97_c3_1523_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l93_c3_cfb0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l85_c7_2701_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_iffalse := VAR_t8_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l96_c7_2fa9] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_cond;
     tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue;
     tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output := tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l90_c7_7d27] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l99_c42_fe5d] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_left;
     BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_return_output := BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;

     -- t8_MUX[uxn_opcodes_h_l85_c7_2701] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l85_c7_2701_cond <= VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_cond;
     t8_MUX_uxn_opcodes_h_l85_c7_2701_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_iftrue;
     t8_MUX_uxn_opcodes_h_l85_c7_2701_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_return_output := t8_MUX_uxn_opcodes_h_l85_c7_2701_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l85_c7_2701] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l90_c7_7d27] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;

     -- Submodule level 3
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_left := VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_fe5d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l85_c7_2701_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l85_c7_2701_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l90_c7_7d27] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_cond;
     tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue;
     tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_return_output := tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l85_c7_2701] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_return_output;

     -- t8_MUX[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l71_c2_beb1_cond <= VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_cond;
     t8_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue;
     t8_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_return_output := t8_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l85_c7_2701] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l99_c42_bc76] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_left;
     BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_return_output := BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_return_output;

     -- Submodule level 4
     VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_iffalse := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l99_c42_bc76_return_output, 16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l85_c7_2701_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l85_c7_2701_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l85_c7_2701] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l85_c7_2701_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_cond;
     tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iftrue;
     tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_return_output := tmp16_MUX_uxn_opcodes_h_l85_c7_2701_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;

     -- MUX[uxn_opcodes_h_l99_c22_e9ee] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l99_c22_e9ee_cond <= VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_cond;
     MUX_uxn_opcodes_h_l99_c22_e9ee_iftrue <= VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_iftrue;
     MUX_uxn_opcodes_h_l99_c22_e9ee_iffalse <= VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_return_output := MUX_uxn_opcodes_h_l99_c22_e9ee_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;

     -- Submodule level 5
     VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue := VAR_MUX_uxn_opcodes_h_l99_c22_e9ee_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l85_c7_2701_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_cond;
     tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue;
     tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_return_output := tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l96_c7_2fa9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output := result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output;

     -- Submodule level 6
     VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l96_c7_2fa9_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l90_c7_7d27] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_cond;
     result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_return_output := result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;

     -- Submodule level 7
     VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l90_c7_7d27_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l85_c7_2701] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_cond;
     result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_return_output := result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_return_output;

     -- Submodule level 8
     VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l85_c7_2701_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l71_c2_beb1] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_cond;
     result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_return_output := result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_161f_uxn_opcodes_h_l103_l66_DUPLICATE_39ef LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_161f_uxn_opcodes_h_l103_l66_DUPLICATE_39ef_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_161f(
     result,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l71_c2_beb1_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l71_c2_beb1_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_161f_uxn_opcodes_h_l103_l66_DUPLICATE_39ef_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_161f_uxn_opcodes_h_l103_l66_DUPLICATE_39ef_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp16 <= REG_COMB_tmp16;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
