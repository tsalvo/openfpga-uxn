-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 66
entity jsr_0CLK_4f993427 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr_0CLK_4f993427;
architecture arch of jsr_0CLK_4f993427 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l712_c6_212b]
signal BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l712_c1_1b91]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l712_c2_f53b]
signal t8_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l712_c2_f53b]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l712_c2_f53b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l712_c2_f53b]
signal result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l712_c2_f53b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l712_c2_f53b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l712_c2_f53b]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l712_c2_f53b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l712_c2_f53b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l712_c2_f53b]
signal result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l713_c3_c418[uxn_opcodes_h_l713_c3_c418]
signal printf_uxn_opcodes_h_l713_c3_c418_uxn_opcodes_h_l713_c3_c418_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l717_c11_41ec]
signal BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l717_c7_ade8]
signal t8_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l717_c7_ade8]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l717_c7_ade8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l717_c7_ade8]
signal result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l717_c7_ade8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l717_c7_ade8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l717_c7_ade8]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l717_c7_ade8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l717_c7_ade8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l717_c7_ade8]
signal result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l720_c11_4889]
signal BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l720_c7_36eb]
signal t8_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l720_c7_36eb]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l720_c7_36eb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l720_c7_36eb]
signal result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l720_c7_36eb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l720_c7_36eb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l720_c7_36eb]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l720_c7_36eb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l720_c7_36eb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l720_c7_36eb]
signal result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l723_c30_ce85]
signal sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l725_c11_5a2f]
signal BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l725_c7_8957]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l725_c7_8957]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l725_c7_8957]
signal result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l725_c7_8957]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l725_c7_8957]
signal result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l725_c7_8957]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l725_c7_8957]
signal result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l725_c7_8957]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l725_c7_8957]
signal result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l732_c11_97db]
signal BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l732_c7_3209]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l732_c7_3209]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l732_c7_3209]
signal result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(15 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l732_c7_3209]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l732_c7_3209]
signal result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l732_c7_3209]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l732_c7_3209]
signal result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l732_c7_3209]
signal result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(7 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l735_c31_0bf7]
signal CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l737_c22_8e34]
signal BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l739_c11_09ef]
signal BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l739_c7_835f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l739_c7_835f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l739_c7_835f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l739_c7_835f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_c785( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.is_stack_write := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b
BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_left,
BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_right,
BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_return_output);

-- t8_MUX_uxn_opcodes_h_l712_c2_f53b
t8_MUX_uxn_opcodes_h_l712_c2_f53b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l712_c2_f53b_cond,
t8_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue,
t8_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse,
t8_MUX_uxn_opcodes_h_l712_c2_f53b_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b
result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b
result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b
result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond,
result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b
result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b
result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b
result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b
result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond,
result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output);

-- printf_uxn_opcodes_h_l713_c3_c418_uxn_opcodes_h_l713_c3_c418
printf_uxn_opcodes_h_l713_c3_c418_uxn_opcodes_h_l713_c3_c418 : entity work.printf_uxn_opcodes_h_l713_c3_c418_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l713_c3_c418_uxn_opcodes_h_l713_c3_c418_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec
BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_left,
BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_right,
BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output);

-- t8_MUX_uxn_opcodes_h_l717_c7_ade8
t8_MUX_uxn_opcodes_h_l717_c7_ade8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l717_c7_ade8_cond,
t8_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue,
t8_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse,
t8_MUX_uxn_opcodes_h_l717_c7_ade8_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8
result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8
result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8
result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond,
result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8
result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8
result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8
result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8
result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond,
result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889
BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_left,
BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_right,
BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output);

-- t8_MUX_uxn_opcodes_h_l720_c7_36eb
t8_MUX_uxn_opcodes_h_l720_c7_36eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l720_c7_36eb_cond,
t8_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue,
t8_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse,
t8_MUX_uxn_opcodes_h_l720_c7_36eb_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb
result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb
result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb
result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond,
result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb
result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb
result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb
result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb
result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond,
result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output);

-- sp_relative_shift_uxn_opcodes_h_l723_c30_ce85
sp_relative_shift_uxn_opcodes_h_l723_c30_ce85 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_ins,
sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_x,
sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_y,
sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f
BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_left,
BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_right,
BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957
result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957
result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957
result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_cond,
result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957
result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957
result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957
result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957
result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_cond,
result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db
BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_left,
BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_right,
BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209
result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209
result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209
result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_cond,
result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209
result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209
result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209
result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_cond,
result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output);

-- CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7
CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_x,
CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34
BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_left,
BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_right,
BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef
BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_left,
BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_right,
BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f
result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f
result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f
result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_return_output,
 t8_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output,
 t8_MUX_uxn_opcodes_h_l717_c7_ade8_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output,
 t8_MUX_uxn_opcodes_h_l720_c7_36eb_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output,
 sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output,
 CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l714_c3_11d6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l713_c3_c418_uxn_opcodes_h_l713_c3_c418_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l718_c3_7f96 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l729_c3_da0c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l727_c3_43ce : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l730_c21_cfb6_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l737_c3_fd94 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l734_c3_9f97 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l735_c21_bb9e_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l737_c27_eb29_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l712_l739_l725_l720_DUPLICATE_a456_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l725_l717_l732_DUPLICATE_eece_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l717_l712_l732_l725_l720_DUPLICATE_bc13_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_da82_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_f7cb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l712_l725_l717_DUPLICATE_f830_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l712_l717_l732_l720_DUPLICATE_73cd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l739_l732_l725_l720_DUPLICATE_e5c7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l732_l720_DUPLICATE_8e5a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c785_uxn_opcodes_h_l746_l708_DUPLICATE_a48d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l714_c3_11d6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l714_c3_11d6;
     VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l729_c3_da0c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l729_c3_da0c;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iffalse := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l734_c3_9f97 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l734_c3_9f97;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_right := to_unsigned(2, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l718_c3_7f96 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l718_c3_7f96;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l727_c3_43ce := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l727_c3_43ce;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse := t8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l732_l720_DUPLICATE_8e5a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l732_l720_DUPLICATE_8e5a_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l717_l712_l732_l725_l720_DUPLICATE_bc13 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l717_l712_l732_l725_l720_DUPLICATE_bc13_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l739_l732_l725_l720_DUPLICATE_e5c7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l739_l732_l725_l720_DUPLICATE_e5c7_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_da82 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_da82_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l725_c11_5a2f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_left;
     BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output := BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l712_l725_l717_DUPLICATE_f830 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l712_l725_l717_DUPLICATE_f830_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l723_c30_ce85] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_ins;
     sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_x <= VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_x;
     sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_y <= VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_return_output := sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l737_c27_eb29] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l737_c27_eb29_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l725_l717_l732_DUPLICATE_eece LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l725_l717_l732_DUPLICATE_eece_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l712_c6_212b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_left;
     BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output := BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_f7cb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_f7cb_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l732_c11_97db] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_left;
     BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output := BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l712_l717_l732_l720_DUPLICATE_73cd LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l712_l717_l732_l720_DUPLICATE_73cd_return_output := result.u8_value;

     -- CONST_SR_8[uxn_opcodes_h_l735_c31_0bf7] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_x <= VAR_CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_return_output := CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l712_l739_l725_l720_DUPLICATE_a456 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l712_l739_l725_l720_DUPLICATE_a456_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l720_c11_4889] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_left;
     BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output := BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l717_c11_41ec] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_left;
     BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output := BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l730_c21_cfb6] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l730_c21_cfb6_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- BIN_OP_EQ[uxn_opcodes_h_l739_c11_09ef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_left;
     BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_return_output := BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l712_c6_212b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l717_c11_41ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l720_c11_4889_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l725_c11_5a2f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l732_c11_97db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l739_c11_09ef_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l737_c27_eb29_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l730_c21_cfb6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l712_l725_l717_DUPLICATE_f830_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l712_l725_l717_DUPLICATE_f830_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l712_l725_l717_DUPLICATE_f830_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l717_l712_l732_l725_l720_DUPLICATE_bc13_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l717_l712_l732_l725_l720_DUPLICATE_bc13_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l717_l712_l732_l725_l720_DUPLICATE_bc13_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l717_l712_l732_l725_l720_DUPLICATE_bc13_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l717_l712_l732_l725_l720_DUPLICATE_bc13_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l739_l732_l725_l720_DUPLICATE_e5c7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l739_l732_l725_l720_DUPLICATE_e5c7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l739_l732_l725_l720_DUPLICATE_e5c7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l739_l732_l725_l720_DUPLICATE_e5c7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l717_l739_l732_l725_l720_DUPLICATE_e5c7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l712_l739_l725_l720_DUPLICATE_a456_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l712_l739_l725_l720_DUPLICATE_a456_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l712_l739_l725_l720_DUPLICATE_a456_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l712_l739_l725_l720_DUPLICATE_a456_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l717_l712_l739_l725_l720_DUPLICATE_a456_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l725_l717_l732_DUPLICATE_eece_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l725_l717_l732_DUPLICATE_eece_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l725_l717_l732_DUPLICATE_eece_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l712_l725_l717_l732_DUPLICATE_eece_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_da82_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_da82_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_da82_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_da82_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_da82_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_f7cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_f7cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_f7cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_f7cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l717_l712_l739_l732_l720_DUPLICATE_f7cb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l732_l720_DUPLICATE_8e5a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l732_l720_DUPLICATE_8e5a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l712_l717_l732_l720_DUPLICATE_73cd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l712_l717_l732_l720_DUPLICATE_73cd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l712_l717_l732_l720_DUPLICATE_73cd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l712_l717_l732_l720_DUPLICATE_73cd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l723_c30_ce85_return_output;
     -- CAST_TO_uint8_t[uxn_opcodes_h_l735_c21_bb9e] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l735_c21_bb9e_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l735_c31_0bf7_return_output);

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l732_c7_3209] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l739_c7_835f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l739_c7_835f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l737_c22_8e34] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_left;
     BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_return_output := BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l739_c7_835f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l712_c1_1b91] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l725_c7_8957] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l732_c7_3209] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l739_c7_835f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_return_output;

     -- t8_MUX[uxn_opcodes_h_l720_c7_36eb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l720_c7_36eb_cond <= VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_cond;
     t8_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue;
     t8_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_return_output := t8_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l737_c3_fd94 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l737_c22_8e34_return_output)),16);
     VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l735_c21_bb9e_return_output;
     VAR_printf_uxn_opcodes_h_l713_c3_c418_uxn_opcodes_h_l713_c3_c418_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l712_c1_1b91_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l739_c7_835f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l739_c7_835f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l732_c7_3209_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l739_c7_835f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l739_c7_835f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l732_c7_3209_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue := VAR_result_u16_value_uxn_opcodes_h_l737_c3_fd94;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l732_c7_3209] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_return_output;

     -- t8_MUX[uxn_opcodes_h_l717_c7_ade8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l717_c7_ade8_cond <= VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_cond;
     t8_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue;
     t8_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_return_output := t8_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l720_c7_36eb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l732_c7_3209] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l732_c7_3209] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l725_c7_8957] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l732_c7_3209] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l732_c7_3209] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_cond;
     result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output := result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output;

     -- printf_uxn_opcodes_h_l713_c3_c418[uxn_opcodes_h_l713_c3_c418] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l713_c3_c418_uxn_opcodes_h_l713_c3_c418_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l713_c3_c418_uxn_opcodes_h_l713_c3_c418_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l732_c7_3209] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_cond;
     result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output := result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l725_c7_8957] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l732_c7_3209_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l732_c7_3209_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l725_c7_8957_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l732_c7_3209_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l732_c7_3209_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l725_c7_8957_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l732_c7_3209_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l725_c7_8957] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l725_c7_8957] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_cond;
     result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output := result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l725_c7_8957] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_cond;
     result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output := result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l717_c7_ade8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l725_c7_8957] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l720_c7_36eb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l725_c7_8957] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l725_c7_8957] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_return_output;

     -- t8_MUX[uxn_opcodes_h_l712_c2_f53b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l712_c2_f53b_cond <= VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_cond;
     t8_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue;
     t8_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_return_output := t8_MUX_uxn_opcodes_h_l712_c2_f53b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l720_c7_36eb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l725_c7_8957_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l725_c7_8957_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l725_c7_8957_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l725_c7_8957_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l725_c7_8957_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l712_c2_f53b_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l720_c7_36eb] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond;
     result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output := result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l720_c7_36eb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l717_c7_ade8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l720_c7_36eb] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l717_c7_ade8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l720_c7_36eb] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l712_c2_f53b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l720_c7_36eb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l720_c7_36eb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output := result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l720_c7_36eb_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l717_c7_ade8] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l717_c7_ade8] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l712_c2_f53b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l717_c7_ade8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l712_c2_f53b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l717_c7_ade8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l717_c7_ade8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output := result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l717_c7_ade8] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_cond;
     result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output := result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l717_c7_ade8_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l712_c2_f53b] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l712_c2_f53b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output := result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l712_c2_f53b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output := result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l712_c2_f53b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l712_c2_f53b] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l712_c2_f53b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c785_uxn_opcodes_h_l746_l708_DUPLICATE_a48d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c785_uxn_opcodes_h_l746_l708_DUPLICATE_a48d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c785(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l712_c2_f53b_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l712_c2_f53b_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c785_uxn_opcodes_h_l746_l708_DUPLICATE_a48d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c785_uxn_opcodes_h_l746_l708_DUPLICATE_a48d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
