-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity ldz_0CLK_f74745d5 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_f74745d5;
architecture arch of ldz_0CLK_f74745d5 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1361_c6_f0f2]
signal BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1361_c1_f2ea]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1361_c2_2294]
signal t8_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1361_c2_2294]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1361_c2_2294]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1361_c2_2294]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1361_c2_2294]
signal result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1361_c2_2294]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1361_c2_2294]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1361_c2_2294]
signal result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(15 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1361_c2_2294]
signal tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1362_c3_c9cc[uxn_opcodes_h_l1362_c3_c9cc]
signal printf_uxn_opcodes_h_l1362_c3_c9cc_uxn_opcodes_h_l1362_c3_c9cc_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1366_c11_6c5c]
signal BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1366_c7_a8d3]
signal t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1366_c7_a8d3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1366_c7_a8d3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1366_c7_a8d3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1366_c7_a8d3]
signal result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1366_c7_a8d3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1366_c7_a8d3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1366_c7_a8d3]
signal result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(15 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1366_c7_a8d3]
signal tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1369_c11_cb85]
signal BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1369_c7_971b]
signal t8_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1369_c7_971b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1369_c7_971b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1369_c7_971b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1369_c7_971b]
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1369_c7_971b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1369_c7_971b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1369_c7_971b]
signal result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(15 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1369_c7_971b]
signal tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1372_c30_7539]
signal sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1375_c11_8f6e]
signal BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1375_c7_a8fd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1375_c7_a8fd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1375_c7_a8fd]
signal result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1375_c7_a8fd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1375_c7_a8fd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1375_c7_a8fd]
signal tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1378_c11_c6cd]
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1378_c7_1d47]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c7_1d47]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c7_1d47]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1378_c7_1d47]
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1378_c7_1d47]
signal tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1384_c11_d42b]
signal BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1384_c7_116b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1384_c7_116b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_ff87( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;
      base.u16_value := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2
BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_left,
BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_right,
BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_return_output);

-- t8_MUX_uxn_opcodes_h_l1361_c2_2294
t8_MUX_uxn_opcodes_h_l1361_c2_2294 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1361_c2_2294_cond,
t8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue,
t8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse,
t8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294
result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294
result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294
result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond,
result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294
result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294
result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294
result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond,
result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1361_c2_2294
tmp8_MUX_uxn_opcodes_h_l1361_c2_2294 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_cond,
tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue,
tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse,
tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output);

-- printf_uxn_opcodes_h_l1362_c3_c9cc_uxn_opcodes_h_l1362_c3_c9cc
printf_uxn_opcodes_h_l1362_c3_c9cc_uxn_opcodes_h_l1362_c3_c9cc : entity work.printf_uxn_opcodes_h_l1362_c3_c9cc_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1362_c3_c9cc_uxn_opcodes_h_l1362_c3_c9cc_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c
BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_left,
BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_right,
BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output);

-- t8_MUX_uxn_opcodes_h_l1366_c7_a8d3
t8_MUX_uxn_opcodes_h_l1366_c7_a8d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond,
t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue,
t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse,
t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3
result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3
result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3
result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3
result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3
result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond,
result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3
tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond,
tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue,
tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse,
tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85
BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_left,
BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_right,
BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output);

-- t8_MUX_uxn_opcodes_h_l1369_c7_971b
t8_MUX_uxn_opcodes_h_l1369_c7_971b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1369_c7_971b_cond,
t8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue,
t8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse,
t8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b
result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b
result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b
result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond,
result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1369_c7_971b
tmp8_MUX_uxn_opcodes_h_l1369_c7_971b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_cond,
tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue,
tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse,
tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1372_c30_7539
sp_relative_shift_uxn_opcodes_h_l1372_c30_7539 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_ins,
sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_x,
sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_y,
sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e
BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_left,
BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_right,
BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd
result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd
result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond,
result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd
result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd
result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd
tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond,
tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue,
tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse,
tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_left,
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_right,
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47
result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_cond,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47
tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_cond,
tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue,
tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse,
tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b
BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_left,
BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_right,
BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b
result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b
result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_return_output,
 t8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
 tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output,
 t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output,
 tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output,
 t8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output,
 tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output,
 sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output,
 tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output,
 tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1363_c3_83f4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1362_c3_c9cc_uxn_opcodes_h_l1362_c3_c9cc_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1367_c3_44d1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1373_c22_49fa_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_9c06 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1366_l1361_l1384_l1375_l1369_DUPLICATE_d760_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_f13f_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1366_l1361_l1378_l1375_l1369_DUPLICATE_f7b5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1361_l1375_l1366_DUPLICATE_914d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_d5b7_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1366_l1384_l1378_l1375_l1369_DUPLICATE_0ad7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1375_l1378_l1369_DUPLICATE_a048_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ff87_uxn_opcodes_h_l1389_l1357_DUPLICATE_94f9_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_9c06 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_9c06;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1363_c3_83f4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1363_c3_83f4;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1367_c3_44d1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1367_c3_44d1;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_right := to_unsigned(5, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1361_c6_f0f2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1378_c11_c6cd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_left;
     BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_return_output := BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_f13f LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_f13f_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1375_c11_8f6e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1366_l1361_l1384_l1375_l1369_DUPLICATE_d760 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1366_l1361_l1384_l1375_l1369_DUPLICATE_d760_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1384_c11_d42b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1372_c30_7539] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_ins;
     sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_x;
     sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_return_output := sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1361_l1375_l1366_DUPLICATE_914d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1361_l1375_l1366_DUPLICATE_914d_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1375_l1378_l1369_DUPLICATE_a048 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1375_l1378_l1369_DUPLICATE_a048_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1369_c11_cb85] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_left;
     BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output := BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_d5b7 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_d5b7_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1366_l1384_l1378_l1375_l1369_DUPLICATE_0ad7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1366_l1384_l1378_l1375_l1369_DUPLICATE_0ad7_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1366_c11_6c5c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1366_l1361_l1378_l1375_l1369_DUPLICATE_f7b5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1366_l1361_l1378_l1375_l1369_DUPLICATE_f7b5_return_output := result.u8_value;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1373_c22_49fa] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1373_c22_49fa_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1361_c6_f0f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1366_c11_6c5c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_cb85_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1375_c11_8f6e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_c6cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1384_c11_d42b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1373_c22_49fa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_f13f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_f13f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_f13f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_d5b7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_d5b7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1361_l1366_l1369_DUPLICATE_d5b7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1366_l1384_l1378_l1375_l1369_DUPLICATE_0ad7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1366_l1384_l1378_l1375_l1369_DUPLICATE_0ad7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1366_l1384_l1378_l1375_l1369_DUPLICATE_0ad7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1366_l1384_l1378_l1375_l1369_DUPLICATE_0ad7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1366_l1384_l1378_l1375_l1369_DUPLICATE_0ad7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1361_l1375_l1366_DUPLICATE_914d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1361_l1375_l1366_DUPLICATE_914d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1361_l1375_l1366_DUPLICATE_914d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1366_l1361_l1384_l1375_l1369_DUPLICATE_d760_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1366_l1361_l1384_l1375_l1369_DUPLICATE_d760_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1366_l1361_l1384_l1375_l1369_DUPLICATE_d760_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1366_l1361_l1384_l1375_l1369_DUPLICATE_d760_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1366_l1361_l1384_l1375_l1369_DUPLICATE_d760_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1375_l1378_l1369_DUPLICATE_a048_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1375_l1378_l1369_DUPLICATE_a048_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1375_l1378_l1369_DUPLICATE_a048_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1366_l1361_l1378_l1375_l1369_DUPLICATE_f7b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1366_l1361_l1378_l1375_l1369_DUPLICATE_f7b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1366_l1361_l1378_l1375_l1369_DUPLICATE_f7b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1366_l1361_l1378_l1375_l1369_DUPLICATE_f7b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1366_l1361_l1378_l1375_l1369_DUPLICATE_f7b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1372_c30_7539_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1375_c7_a8fd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1384_c7_116b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1369_c7_971b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output := result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1378_c7_1d47] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_cond;
     tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output := tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1378_c7_1d47] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output := result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1369_c7_971b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1369_c7_971b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1369_c7_971b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_cond;
     t8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue;
     t8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output := t8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1361_c1_f2ea] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c7_1d47] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1384_c7_116b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1362_c3_c9cc_uxn_opcodes_h_l1362_c3_c9cc_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1361_c1_f2ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1384_c7_116b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1384_c7_116b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output;
     -- printf_uxn_opcodes_h_l1362_c3_c9cc[uxn_opcodes_h_l1362_c3_c9cc] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1362_c3_c9cc_uxn_opcodes_h_l1362_c3_c9cc_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1362_c3_c9cc_uxn_opcodes_h_l1362_c3_c9cc_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1375_c7_a8fd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1375_c7_a8fd] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond;
     tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output := tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1369_c7_971b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1366_c7_a8d3] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output := result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;

     -- t8_MUX[uxn_opcodes_h_l1366_c7_a8d3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond <= VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond;
     t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue;
     t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output := t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1375_c7_a8fd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output := result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1366_c7_a8d3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c7_1d47] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1378_c7_1d47] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c7_1d47_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1369_c7_971b] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_cond;
     tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output := tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1361_c2_2294] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1361_c2_2294_cond <= VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_cond;
     t8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue;
     t8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output := t8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1361_c2_2294] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1369_c7_971b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1375_c7_a8fd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1369_c7_971b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1361_c2_2294] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output := result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1375_c7_a8fd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1366_c7_a8d3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1375_c7_a8fd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1366_c7_a8d3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1366_c7_a8d3] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond;
     tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output := tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1369_c7_971b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1366_c7_a8d3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1361_c2_2294] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1369_c7_971b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_971b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1361_c2_2294] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1361_c2_2294] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output := result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1361_c2_2294] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_cond;
     tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output := tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1366_c7_a8d3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1366_c7_a8d3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1366_c7_a8d3_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1361_c2_2294_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1361_c2_2294] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1361_c2_2294] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_ff87_uxn_opcodes_h_l1389_l1357_DUPLICATE_94f9 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ff87_uxn_opcodes_h_l1389_l1357_DUPLICATE_94f9_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_ff87(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1361_c2_2294_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1361_c2_2294_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ff87_uxn_opcodes_h_l1389_l1357_DUPLICATE_94f9_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ff87_uxn_opcodes_h_l1389_l1357_DUPLICATE_94f9_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
