-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity lit2_0CLK_4c8178ef is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lit2_0CLK_4c8178ef;
architecture arch of lit2_0CLK_4c8178ef is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l222_c6_240a]
signal BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l222_c2_e06f]
signal result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l222_c2_e06f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l222_c2_e06f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l222_c2_e06f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l222_c2_e06f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l222_c2_e06f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l222_c2_e06f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l222_c2_e06f]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l222_c2_e06f]
signal tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l231_c11_3cb4]
signal BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l231_c7_20f9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l231_c7_20f9]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l231_c7_20f9]
signal result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l231_c7_20f9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l231_c7_20f9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l231_c7_20f9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l231_c7_20f9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(3 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l231_c7_20f9]
signal tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l233_c22_285e]
signal BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l235_c11_df7d]
signal BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l235_c7_796f]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l235_c7_796f]
signal result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l235_c7_796f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l235_c7_796f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l235_c7_796f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l235_c7_796f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(3 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l235_c7_796f]
signal tmp16_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l237_c3_42f2]
signal CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l239_c22_0a0a]
signal BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_right : unsigned(1 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l241_c11_8334]
signal BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l241_c7_cb50]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l241_c7_cb50]
signal result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l241_c7_cb50]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l241_c7_cb50]
signal result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l241_c7_cb50]
signal result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l241_c7_cb50]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(3 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l241_c7_cb50]
signal tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l242_c3_baee]
signal BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l249_c11_1ba6]
signal BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l249_c7_dddb]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l249_c7_dddb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l249_c7_dddb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_41b6( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_sp_shift := ref_toks_7;
      base.is_stack_operation_16bit := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a
BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_left,
BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_right,
BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f
result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_cond,
result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f
result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f
result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f
result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f
result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f
result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_return_output);

-- tmp16_MUX_uxn_opcodes_h_l222_c2_e06f
tmp16_MUX_uxn_opcodes_h_l222_c2_e06f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_cond,
tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue,
tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse,
tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4
BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_left,
BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_right,
BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9
result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9
result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_cond,
result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9
result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9
result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9
result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_return_output);

-- tmp16_MUX_uxn_opcodes_h_l231_c7_20f9
tmp16_MUX_uxn_opcodes_h_l231_c7_20f9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_cond,
tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue,
tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse,
tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e
BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_left,
BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_right,
BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d
BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_left,
BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_right,
BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f
result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_cond,
result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f
result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f
result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f
result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_return_output);

-- tmp16_MUX_uxn_opcodes_h_l235_c7_796f
tmp16_MUX_uxn_opcodes_h_l235_c7_796f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l235_c7_796f_cond,
tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iftrue,
tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iffalse,
tmp16_MUX_uxn_opcodes_h_l235_c7_796f_return_output);

-- CONST_SL_8_uxn_opcodes_h_l237_c3_42f2
CONST_SL_8_uxn_opcodes_h_l237_c3_42f2 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_x,
CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a
BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a : entity work.BIN_OP_PLUS_uint16_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_left,
BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_right,
BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334
BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_left,
BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_right,
BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50
result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_cond,
result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50
result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50
result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50
result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_return_output);

-- tmp16_MUX_uxn_opcodes_h_l241_c7_cb50
tmp16_MUX_uxn_opcodes_h_l241_c7_cb50 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_cond,
tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue,
tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse,
tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l242_c3_baee
BIN_OP_OR_uxn_opcodes_h_l242_c3_baee : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_left,
BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_right,
BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6
BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_left,
BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_right,
BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb
result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb
result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_ram_read,
 -- Registers
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
 tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_return_output,
 tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_return_output,
 tmp16_MUX_uxn_opcodes_h_l235_c7_796f_return_output,
 CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_return_output,
 tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_return_output,
 BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l227_c3_c874 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l222_c2_e06f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l231_c7_20f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l233_c3_48b5 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l239_c3_014e : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l241_c7_cb50_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l245_c3_846c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l222_l241_l231_DUPLICATE_7e6c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_c42b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l235_l222_l241_l231_DUPLICATE_be2f_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_929a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l235_l241_l231_l249_DUPLICATE_792c_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l236_l242_DUPLICATE_c719_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_41b6_uxn_opcodes_h_l255_l217_DUPLICATE_2e89_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_right := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l227_c3_c874 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l227_c3_c874;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_right := to_unsigned(2, 2);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l245_c3_846c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l245_c3_846c;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_left := VAR_pc;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_left := VAR_pc;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_left := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse := tmp16;
     -- BIN_OP_EQ[uxn_opcodes_h_l249_c11_1ba6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_left;
     BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_return_output := BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l235_l222_l241_l231_DUPLICATE_be2f LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l235_l222_l241_l231_DUPLICATE_be2f_return_output := result.stack_address_sp_offset;

     -- BIN_OP_PLUS[uxn_opcodes_h_l239_c22_0a0a] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_left;
     BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_return_output := BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l222_c6_240a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_left;
     BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output := BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l235_l241_l231_l249_DUPLICATE_792c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l235_l241_l231_l249_DUPLICATE_792c_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l231_c11_3cb4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_left;
     BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output := BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l235_c11_df7d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_left;
     BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output := BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output;

     -- result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d[uxn_opcodes_h_l231_c7_20f9] LATENCY=0
     VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l231_c7_20f9_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_929a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_929a_return_output := result.is_stack_operation_16bit;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l222_c2_e06f] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l222_c2_e06f_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_c42b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_c42b_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l222_l241_l231_DUPLICATE_7e6c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l222_l241_l231_DUPLICATE_7e6c_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l241_c11_8334] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_left;
     BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output := BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l233_c22_285e] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_left;
     BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_return_output := BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l236_l242_DUPLICATE_c719 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l236_l242_DUPLICATE_c719_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_ram_read);

     -- result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d[uxn_opcodes_h_l241_c7_cb50] LATENCY=0
     VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l241_c7_cb50_return_output := result.u16_value;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l222_c6_240a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l231_c11_3cb4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l235_c11_df7d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l241_c11_8334_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l249_c11_1ba6_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l233_c3_48b5 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l233_c22_285e_return_output, 16);
     VAR_result_u16_value_uxn_opcodes_h_l239_c3_014e := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l239_c22_0a0a_return_output, 16);
     VAR_BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l236_l242_DUPLICATE_c719_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l236_l242_DUPLICATE_c719_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l235_l241_l231_l249_DUPLICATE_792c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l235_l241_l231_l249_DUPLICATE_792c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l235_l241_l231_l249_DUPLICATE_792c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l235_l241_l231_l249_DUPLICATE_792c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l222_l241_l231_DUPLICATE_7e6c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l222_l241_l231_DUPLICATE_7e6c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l222_l241_l231_DUPLICATE_7e6c_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_929a_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_929a_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_929a_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_929a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_c42b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_c42b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_c42b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l235_l222_l231_l249_DUPLICATE_c42b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l235_l222_l241_l231_DUPLICATE_be2f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l235_l222_l241_l231_DUPLICATE_be2f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l235_l222_l241_l231_DUPLICATE_be2f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l235_l222_l241_l231_DUPLICATE_be2f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse := VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l231_c7_20f9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l222_c2_e06f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse := VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l241_c7_cb50_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue := VAR_result_u16_value_uxn_opcodes_h_l233_c3_48b5;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iftrue := VAR_result_u16_value_uxn_opcodes_h_l239_c3_014e;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l231_c7_20f9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l249_c7_dddb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l237_c3_42f2] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_x <= VAR_CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_return_output := CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l241_c7_cb50] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l249_c7_dddb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l241_c7_cb50] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l242_c3_baee] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_left;
     BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_return_output := BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l249_c7_dddb] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l222_c2_e06f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output;

     -- Submodule level 2
     VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l242_c3_baee_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l237_c3_42f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l249_c7_dddb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l249_c7_dddb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l249_c7_dddb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l222_c2_e06f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l235_c7_796f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l241_c7_cb50] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l241_c7_cb50] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_cond;
     result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_return_output := result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l241_c7_cb50] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l235_c7_796f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l241_c7_cb50] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l241_c7_cb50] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_cond;
     tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iftrue;
     tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_return_output := tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l235_c7_796f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l235_c7_796f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l241_c7_cb50_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l235_c7_796f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l235_c7_796f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l235_c7_796f] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l235_c7_796f_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_cond;
     tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iftrue;
     tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_return_output := tmp16_MUX_uxn_opcodes_h_l235_c7_796f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l231_c7_20f9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l235_c7_796f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_return_output := result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l231_c7_20f9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l235_c7_796f] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l235_c7_796f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l235_c7_796f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l235_c7_796f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l235_c7_796f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l235_c7_796f_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l222_c2_e06f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l231_c7_20f9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l231_c7_20f9] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l222_c2_e06f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l231_c7_20f9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_return_output := result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l231_c7_20f9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l231_c7_20f9] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_cond;
     tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iftrue;
     tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_return_output := tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l231_c7_20f9_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l222_c2_e06f] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_cond;
     tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue;
     tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_return_output := tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l222_c2_e06f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l222_c2_e06f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_return_output := result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l222_c2_e06f] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l222_c2_e06f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_return_output;

     -- Submodule level 6
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l222_c2_e06f_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_41b6_uxn_opcodes_h_l255_l217_DUPLICATE_2e89 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_41b6_uxn_opcodes_h_l255_l217_DUPLICATE_2e89_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_41b6(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l222_c2_e06f_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l222_c2_e06f_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_41b6_uxn_opcodes_h_l255_l217_DUPLICATE_2e89_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_41b6_uxn_opcodes_h_l255_l217_DUPLICATE_2e89_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
