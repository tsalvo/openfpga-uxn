-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 42
entity sth_0CLK_61914e8d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_61914e8d;
architecture arch of sth_0CLK_61914e8d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2540_c6_e44b]
signal BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2540_c2_93b6]
signal t8_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2540_c2_93b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2540_c2_93b6]
signal result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2540_c2_93b6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2540_c2_93b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2540_c2_93b6]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2540_c2_93b6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2540_c2_93b6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2545_c11_62c3]
signal BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2545_c7_c464]
signal t8_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2545_c7_c464]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2545_c7_c464]
signal result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2545_c7_c464]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2545_c7_c464]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2545_c7_c464]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2545_c7_c464]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2545_c7_c464]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2548_c11_5eab]
signal BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2548_c7_d44c]
signal t8_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2548_c7_d44c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2548_c7_d44c]
signal result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2548_c7_d44c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2548_c7_d44c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2548_c7_d44c]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2548_c7_d44c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2548_c7_d44c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2551_c30_f1b7]
signal sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2553_c11_1d40]
signal BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2553_c7_cf5c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2553_c7_cf5c]
signal result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2553_c7_cf5c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2553_c7_cf5c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2553_c7_cf5c]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2553_c7_cf5c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2553_c7_cf5c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2560_c11_c7cf]
signal BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2560_c7_0b4a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2560_c7_0b4a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2560_c7_0b4a]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2560_c7_0b4a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_4605( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_sp_shift := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b
BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_left,
BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_right,
BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output);

-- t8_MUX_uxn_opcodes_h_l2540_c2_93b6
t8_MUX_uxn_opcodes_h_l2540_c2_93b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2540_c2_93b6_cond,
t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue,
t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse,
t8_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6
result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6
result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6
result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6
result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3
BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_left,
BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_right,
BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output);

-- t8_MUX_uxn_opcodes_h_l2545_c7_c464
t8_MUX_uxn_opcodes_h_l2545_c7_c464 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2545_c7_c464_cond,
t8_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue,
t8_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse,
t8_MUX_uxn_opcodes_h_l2545_c7_c464_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464
result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_cond,
result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464
result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464
result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464
result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464
result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab
BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_left,
BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_right,
BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output);

-- t8_MUX_uxn_opcodes_h_l2548_c7_d44c
t8_MUX_uxn_opcodes_h_l2548_c7_d44c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2548_c7_d44c_cond,
t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue,
t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse,
t8_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c
result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c
result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c
result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c
result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7
sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_ins,
sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_x,
sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_y,
sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40
BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_left,
BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_right,
BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c
result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c
result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c
result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c
result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf
BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_left,
BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_right,
BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a
result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a
result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a
result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output,
 t8_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output,
 t8_MUX_uxn_opcodes_h_l2545_c7_c464_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output,
 t8_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output,
 sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2542_c3_29dd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2546_c3_98a0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2557_c3_ec14 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2555_c3_0530 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2553_l2545_l2548_l2540_DUPLICATE_ebdf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_fdec_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_c99d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2553_l2545_l2540_DUPLICATE_9407_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2540_DUPLICATE_97b7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2548_DUPLICATE_4955_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2553_l2548_DUPLICATE_2843_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4605_uxn_opcodes_h_l2536_l2567_DUPLICATE_68ff_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2557_c3_ec14 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2557_c3_ec14;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2555_c3_0530 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2555_c3_0530;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_right := to_unsigned(4, 3);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2542_c3_29dd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2542_c3_29dd;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2546_c3_98a0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2546_c3_98a0;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2560_c11_c7cf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_left;
     BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_return_output := BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2553_l2548_DUPLICATE_2843 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2553_l2548_DUPLICATE_2843_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2548_DUPLICATE_4955 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2548_DUPLICATE_4955_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2545_c11_62c3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_c99d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_c99d_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2540_c6_e44b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2553_c11_1d40] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_left;
     BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output := BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2553_l2545_l2548_l2540_DUPLICATE_ebdf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2553_l2545_l2548_l2540_DUPLICATE_ebdf_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2553_l2545_l2540_DUPLICATE_9407 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2553_l2545_l2540_DUPLICATE_9407_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2540_DUPLICATE_97b7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2540_DUPLICATE_97b7_return_output := result.is_sp_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2551_c30_f1b7] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_ins;
     sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_x;
     sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_return_output := sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_fdec LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_fdec_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2548_c11_5eab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_left;
     BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output := BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2540_c6_e44b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2545_c11_62c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2548_c11_5eab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2553_c11_1d40_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2560_c11_c7cf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2553_l2545_l2540_DUPLICATE_9407_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2553_l2545_l2540_DUPLICATE_9407_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2553_l2545_l2540_DUPLICATE_9407_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2548_DUPLICATE_4955_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2548_DUPLICATE_4955_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2548_DUPLICATE_4955_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2548_DUPLICATE_4955_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2540_DUPLICATE_97b7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2540_DUPLICATE_97b7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2540_DUPLICATE_97b7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2553_l2545_l2560_l2540_DUPLICATE_97b7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_c99d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_c99d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_c99d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_c99d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_fdec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_fdec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_fdec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2545_l2560_l2548_l2540_DUPLICATE_fdec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2553_l2548_DUPLICATE_2843_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2553_l2548_DUPLICATE_2843_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2553_l2545_l2548_l2540_DUPLICATE_ebdf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2553_l2545_l2548_l2540_DUPLICATE_ebdf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2553_l2545_l2548_l2540_DUPLICATE_ebdf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2553_l2545_l2548_l2540_DUPLICATE_ebdf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2551_c30_f1b7_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2560_c7_0b4a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2560_c7_0b4a] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2553_c7_cf5c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2560_c7_0b4a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2553_c7_cf5c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2553_c7_cf5c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2560_c7_0b4a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output;

     -- t8_MUX[uxn_opcodes_h_l2548_c7_d44c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2548_c7_d44c_cond <= VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_cond;
     t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue;
     t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output := t8_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2560_c7_0b4a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2553_c7_cf5c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;

     -- t8_MUX[uxn_opcodes_h_l2545_c7_c464] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2545_c7_c464_cond <= VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_cond;
     t8_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue;
     t8_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_return_output := t8_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2548_c7_d44c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2553_c7_cf5c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2553_c7_cf5c] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2548_c7_d44c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2548_c7_d44c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2553_c7_cf5c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2553_c7_cf5c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2548_c7_d44c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2548_c7_d44c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2548_c7_d44c] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;

     -- t8_MUX[uxn_opcodes_h_l2540_c2_93b6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2540_c2_93b6_cond <= VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_cond;
     t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue;
     t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output := t8_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2545_c7_c464] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2548_c7_d44c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2545_c7_c464] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2545_c7_c464] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_return_output := result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2548_c7_d44c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2545_c7_c464] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2545_c7_c464] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2545_c7_c464] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2545_c7_c464] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2540_c2_93b6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2540_c2_93b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2540_c2_93b6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2545_c7_c464_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2540_c2_93b6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2540_c2_93b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2540_c2_93b6] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2540_c2_93b6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4605_uxn_opcodes_h_l2536_l2567_DUPLICATE_68ff LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4605_uxn_opcodes_h_l2536_l2567_DUPLICATE_68ff_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4605(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2540_c2_93b6_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4605_uxn_opcodes_h_l2536_l2567_DUPLICATE_68ff_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4605_uxn_opcodes_h_l2536_l2567_DUPLICATE_68ff_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
