-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity mul_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end mul_0CLK_f62d646e;
architecture arch of mul_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2097_c6_ef8e]
signal BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2097_c1_6886]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2097_c2_3a97]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2097_c2_3a97]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2097_c2_3a97]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2097_c2_3a97]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2097_c2_3a97]
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2097_c2_3a97]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2097_c2_3a97]
signal t8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2097_c2_3a97]
signal n8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2098_c3_6076[uxn_opcodes_h_l2098_c3_6076]
signal printf_uxn_opcodes_h_l2098_c3_6076_uxn_opcodes_h_l2098_c3_6076_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2102_c11_b335]
signal BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2102_c7_1c04]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2102_c7_1c04]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2102_c7_1c04]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2102_c7_1c04]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2102_c7_1c04]
signal result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2102_c7_1c04]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2102_c7_1c04]
signal t8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2102_c7_1c04]
signal n8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2105_c11_938b]
signal BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2105_c7_a663]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2105_c7_a663]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2105_c7_a663]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2105_c7_a663]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2105_c7_a663]
signal result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2105_c7_a663]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2105_c7_a663]
signal t8_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2105_c7_a663]
signal n8_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2109_c11_4219]
signal BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2109_c7_9894]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2109_c7_9894]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2109_c7_9894]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2109_c7_9894]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2109_c7_9894]
signal result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2109_c7_9894]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2109_c7_9894]
signal n8_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2112_c11_2d53]
signal BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2112_c7_f58b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2112_c7_f58b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2112_c7_f58b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2112_c7_f58b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2112_c7_f58b]
signal result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2112_c7_f58b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2112_c7_f58b]
signal n8_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2115_c30_c00a]
signal sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_return_output : signed(3 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l2118_c21_e3de]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2120_c11_df31]
signal BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2120_c7_c62e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2120_c7_c62e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2120_c7_c62e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e
BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_left,
BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_right,
BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97
result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97
result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_cond,
result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output);

-- t8_MUX_uxn_opcodes_h_l2097_c2_3a97
t8_MUX_uxn_opcodes_h_l2097_c2_3a97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond,
t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue,
t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse,
t8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output);

-- n8_MUX_uxn_opcodes_h_l2097_c2_3a97
n8_MUX_uxn_opcodes_h_l2097_c2_3a97 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond,
n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue,
n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse,
n8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output);

-- printf_uxn_opcodes_h_l2098_c3_6076_uxn_opcodes_h_l2098_c3_6076
printf_uxn_opcodes_h_l2098_c3_6076_uxn_opcodes_h_l2098_c3_6076 : entity work.printf_uxn_opcodes_h_l2098_c3_6076_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2098_c3_6076_uxn_opcodes_h_l2098_c3_6076_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335
BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_left,
BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_right,
BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04
result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04
result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04
result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04
result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_cond,
result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04
result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output);

-- t8_MUX_uxn_opcodes_h_l2102_c7_1c04
t8_MUX_uxn_opcodes_h_l2102_c7_1c04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond,
t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue,
t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse,
t8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output);

-- n8_MUX_uxn_opcodes_h_l2102_c7_1c04
n8_MUX_uxn_opcodes_h_l2102_c7_1c04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond,
n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue,
n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse,
n8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b
BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_left,
BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_right,
BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663
result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663
result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663
result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663
result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_cond,
result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663
result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output);

-- t8_MUX_uxn_opcodes_h_l2105_c7_a663
t8_MUX_uxn_opcodes_h_l2105_c7_a663 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2105_c7_a663_cond,
t8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue,
t8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse,
t8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output);

-- n8_MUX_uxn_opcodes_h_l2105_c7_a663
n8_MUX_uxn_opcodes_h_l2105_c7_a663 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2105_c7_a663_cond,
n8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue,
n8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse,
n8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219
BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_left,
BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_right,
BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894
result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894
result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894
result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894
result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_cond,
result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894
result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output);

-- n8_MUX_uxn_opcodes_h_l2109_c7_9894
n8_MUX_uxn_opcodes_h_l2109_c7_9894 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2109_c7_9894_cond,
n8_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue,
n8_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse,
n8_MUX_uxn_opcodes_h_l2109_c7_9894_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53
BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_left,
BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_right,
BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b
result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b
result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b
result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b
result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output);

-- n8_MUX_uxn_opcodes_h_l2112_c7_f58b
n8_MUX_uxn_opcodes_h_l2112_c7_f58b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2112_c7_f58b_cond,
n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue,
n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse,
n8_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a
sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_ins,
sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_x,
sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_y,
sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31
BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_left,
BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_right,
BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e
result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e
result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e
result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
 t8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
 n8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output,
 t8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output,
 n8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output,
 t8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output,
 n8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output,
 n8_MUX_uxn_opcodes_h_l2109_c7_9894_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output,
 n8_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output,
 sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2099_c3_fbf2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2098_c3_6076_uxn_opcodes_h_l2098_c3_6076_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2103_c3_0996 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2107_c3_222b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2110_c3_c78c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2117_c3_adcb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2112_c7_f58b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l2118_c3_6a49 : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_87e8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_6665_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_5db8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_4044_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2102_l2120_l2112_l2109_l2105_DUPLICATE_cf2c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2126_l2093_DUPLICATE_d995_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2110_c3_c78c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2110_c3_c78c;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2117_c3_adcb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2117_c3_adcb;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2099_c3_fbf2 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2099_c3_fbf2;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2103_c3_0996 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2103_c3_0996;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2107_c3_222b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2107_c3_222b;
     VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_left := VAR_phase;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2109_c11_4219] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_left;
     BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output := BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_4044 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_4044_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2097_c6_ef8e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2120_c11_df31] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_left;
     BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_return_output := BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_6665 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_6665_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2112_c11_2d53] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_left;
     BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output := BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2102_l2120_l2112_l2109_l2105_DUPLICATE_cf2c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2102_l2120_l2112_l2109_l2105_DUPLICATE_cf2c_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2102_c11_b335] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_left;
     BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output := BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l2118_c21_e3de] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_5db8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_5db8_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_87e8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_87e8_return_output := result.is_sp_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2112_c7_f58b] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2112_c7_f58b_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l2115_c30_c00a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_ins;
     sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_x;
     sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_return_output := sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2105_c11_938b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c6_ef8e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c11_b335_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2105_c11_938b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2109_c11_4219_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2112_c11_2d53_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2120_c11_df31_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l2118_c3_6a49 := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2118_c21_e3de_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_4044_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_4044_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_4044_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_4044_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_4044_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2102_l2120_l2112_l2109_l2105_DUPLICATE_cf2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2102_l2120_l2112_l2109_l2105_DUPLICATE_cf2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2102_l2120_l2112_l2109_l2105_DUPLICATE_cf2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2102_l2120_l2112_l2109_l2105_DUPLICATE_cf2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2102_l2120_l2112_l2109_l2105_DUPLICATE_cf2c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_87e8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_87e8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_87e8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_87e8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_87e8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_6665_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_6665_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_6665_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_6665_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2102_l2097_l2120_l2109_l2105_DUPLICATE_6665_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_5db8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_5db8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_5db8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_5db8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2102_l2097_l2112_l2109_l2105_DUPLICATE_5db8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2112_c7_f58b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2115_c30_c00a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue := VAR_result_u8_value_uxn_opcodes_h_l2118_c3_6a49;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2112_c7_f58b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2112_c7_f58b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2120_c7_c62e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2120_c7_c62e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2097_c1_6886] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2112_c7_f58b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;

     -- t8_MUX[uxn_opcodes_h_l2105_c7_a663] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2105_c7_a663_cond <= VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_cond;
     t8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue;
     t8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output := t8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2120_c7_c62e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2112_c7_f58b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2112_c7_f58b_cond <= VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_cond;
     n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue;
     n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output := n8_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2098_c3_6076_uxn_opcodes_h_l2098_c3_6076_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2097_c1_6886_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2120_c7_c62e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;
     -- n8_MUX[uxn_opcodes_h_l2109_c7_9894] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2109_c7_9894_cond <= VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_cond;
     n8_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue;
     n8_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_return_output := n8_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2112_c7_f58b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2109_c7_9894] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2109_c7_9894] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_return_output := result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2112_c7_f58b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;

     -- t8_MUX[uxn_opcodes_h_l2102_c7_1c04] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond <= VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond;
     t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue;
     t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output := t8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2112_c7_f58b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2109_c7_9894] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;

     -- printf_uxn_opcodes_h_l2098_c3_6076[uxn_opcodes_h_l2098_c3_6076] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2098_c3_6076_uxn_opcodes_h_l2098_c3_6076_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2098_c3_6076_uxn_opcodes_h_l2098_c3_6076_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2112_c7_f58b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2109_c7_9894] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;

     -- t8_MUX[uxn_opcodes_h_l2097_c2_3a97] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond <= VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond;
     t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue;
     t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output := t8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output;

     -- n8_MUX[uxn_opcodes_h_l2105_c7_a663] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2105_c7_a663_cond <= VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_cond;
     n8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue;
     n8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output := n8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2105_c7_a663] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2105_c7_a663] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_return_output := result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2109_c7_9894] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2109_c7_9894] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2105_c7_a663] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2109_c7_9894_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2102_c7_1c04] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;

     -- n8_MUX[uxn_opcodes_h_l2102_c7_1c04] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond <= VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_cond;
     n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue;
     n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output := n8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2105_c7_a663] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2102_c7_1c04] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2102_c7_1c04] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output := result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2105_c7_a663] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2105_c7_a663] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2105_c7_a663_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2102_c7_1c04] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2097_c2_3a97] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output;

     -- n8_MUX[uxn_opcodes_h_l2097_c2_3a97] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond <= VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_cond;
     n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue;
     n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output := n8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2097_c2_3a97] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output := result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2102_c7_1c04] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2097_c2_3a97] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2102_c7_1c04] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2102_c7_1c04_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2097_c2_3a97] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2097_c2_3a97] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2097_c2_3a97] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2126_l2093_DUPLICATE_d995 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2126_l2093_DUPLICATE_d995_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c2_3a97_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2126_l2093_DUPLICATE_d995_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l2126_l2093_DUPLICATE_d995_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
