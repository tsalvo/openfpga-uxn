-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity ldr_0CLK_a6885b22 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_a6885b22;
architecture arch of ldr_0CLK_a6885b22 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1689_c6_d44a]
signal BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1689_c1_7a1c]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1689_c2_7f74]
signal tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1689_c2_7f74]
signal t8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1689_c2_7f74]
signal result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1689_c2_7f74]
signal result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1689_c2_7f74]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1689_c2_7f74]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1689_c2_7f74]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1689_c2_7f74]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1689_c2_7f74]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(3 downto 0);

-- printf_uxn_opcodes_h_l1690_c3_acb9[uxn_opcodes_h_l1690_c3_acb9]
signal printf_uxn_opcodes_h_l1690_c3_acb9_uxn_opcodes_h_l1690_c3_acb9_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1694_c11_5b6c]
signal BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1694_c7_6df0]
signal tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1694_c7_6df0]
signal t8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1694_c7_6df0]
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1694_c7_6df0]
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1694_c7_6df0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1694_c7_6df0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1694_c7_6df0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1694_c7_6df0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1694_c7_6df0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1697_c11_73bc]
signal BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1697_c7_76b8]
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1697_c7_76b8]
signal t8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1697_c7_76b8]
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1697_c7_76b8]
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1697_c7_76b8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1697_c7_76b8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1697_c7_76b8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1697_c7_76b8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1697_c7_76b8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1700_c30_b49e]
signal sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1701_c22_eddc]
signal BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1703_c11_0dfd]
signal BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1703_c7_e5bb]
signal tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1703_c7_e5bb]
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1703_c7_e5bb]
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1703_c7_e5bb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1703_c7_e5bb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1703_c7_e5bb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1703_c7_e5bb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1705_c22_3c8e]
signal BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1707_c11_464c]
signal BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1707_c7_c931]
signal tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1707_c7_c931]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1707_c7_c931]
signal result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1707_c7_c931]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1707_c7_c931]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1713_c11_2531]
signal BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1713_c7_1319]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1713_c7_1319]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_9969( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.u16_value := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_sp_shift := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a
BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_left,
BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_right,
BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74
tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond,
tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue,
tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse,
tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output);

-- t8_MUX_uxn_opcodes_h_l1689_c2_7f74
t8_MUX_uxn_opcodes_h_l1689_c2_7f74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond,
t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue,
t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse,
t8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74
result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond,
result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74
result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond,
result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74
result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74
result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74
result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74
result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output);

-- printf_uxn_opcodes_h_l1690_c3_acb9_uxn_opcodes_h_l1690_c3_acb9
printf_uxn_opcodes_h_l1690_c3_acb9_uxn_opcodes_h_l1690_c3_acb9 : entity work.printf_uxn_opcodes_h_l1690_c3_acb9_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1690_c3_acb9_uxn_opcodes_h_l1690_c3_acb9_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c
BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_left,
BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_right,
BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0
tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond,
tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue,
tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse,
tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output);

-- t8_MUX_uxn_opcodes_h_l1694_c7_6df0
t8_MUX_uxn_opcodes_h_l1694_c7_6df0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond,
t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue,
t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse,
t8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0
result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0
result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond,
result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_left,
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_right,
BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8
tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond,
tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue,
tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse,
tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output);

-- t8_MUX_uxn_opcodes_h_l1697_c7_76b8
t8_MUX_uxn_opcodes_h_l1697_c7_76b8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond,
t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue,
t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse,
t8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond,
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond,
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e
sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_ins,
sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_x,
sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_y,
sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc
BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_left,
BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_right,
BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_left,
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_right,
BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb
tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond,
tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue,
tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse,
tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond,
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond,
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb
result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb
result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e
BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_left,
BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_right,
BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c
BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_left,
BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_right,
BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1707_c7_c931
tmp8_MUX_uxn_opcodes_h_l1707_c7_c931 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_cond,
tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue,
tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse,
tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931
result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931
result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_cond,
result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931
result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531
BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_left,
BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_right,
BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319
result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319
result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
 t8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output,
 t8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output,
 tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output,
 t8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output,
 sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output,
 tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iffalse : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1691_c3_ae21 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1690_c3_acb9_uxn_opcodes_h_l1690_c3_acb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1695_c3_98d0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1701_c3_ca3e : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1701_c27_048d_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1705_c3_1917 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1705_c27_d911_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1710_c3_8cd2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_9eca_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_075d_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_cb85_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1713_l1703_l1697_l1694_l1689_DUPLICATE_53dc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_cac1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1713_l1707_l1703_l1697_l1694_DUPLICATE_222a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_f825_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9969_uxn_opcodes_h_l1685_l1718_DUPLICATE_3ec6_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1691_c3_ae21 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1691_c3_ae21;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1695_c3_98d0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1695_c3_98d0;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1710_c3_8cd2 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1710_c3_8cd2;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1697_c11_73bc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_left;
     BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output := BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1707_c11_464c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1713_c11_2531] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_left;
     BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_return_output := BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_cb85 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_cb85_return_output := result.sp_relative_shift;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1705_c27_d911] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1705_c27_d911_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_9eca LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_9eca_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1694_c11_5b6c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1713_l1703_l1697_l1694_l1689_DUPLICATE_53dc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1713_l1703_l1697_l1694_l1689_DUPLICATE_53dc_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_f825 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_f825_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1703_c11_0dfd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_left;
     BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output := BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1713_l1707_l1703_l1697_l1694_DUPLICATE_222a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1713_l1707_l1703_l1697_l1694_DUPLICATE_222a_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_cac1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_cac1_return_output := result.is_sp_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1700_c30_b49e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_ins;
     sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_x;
     sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_return_output := sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1701_c27_048d] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1701_c27_048d_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l1689_c6_d44a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_075d LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_075d_return_output := result.u16_value;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1689_c6_d44a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1694_c11_5b6c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1697_c11_73bc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1703_c11_0dfd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1707_c11_464c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1713_c11_2531_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1701_c27_048d_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1705_c27_d911_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_cb85_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_cb85_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1694_l1697_l1689_DUPLICATE_cb85_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_075d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_075d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_075d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1713_l1707_l1703_l1697_l1694_DUPLICATE_222a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1713_l1707_l1703_l1697_l1694_DUPLICATE_222a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1713_l1707_l1703_l1697_l1694_DUPLICATE_222a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1713_l1707_l1703_l1697_l1694_DUPLICATE_222a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1713_l1707_l1703_l1697_l1694_DUPLICATE_222a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_cac1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_cac1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1694_l1689_l1703_DUPLICATE_cac1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1713_l1703_l1697_l1694_l1689_DUPLICATE_53dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1713_l1703_l1697_l1694_l1689_DUPLICATE_53dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1713_l1703_l1697_l1694_l1689_DUPLICATE_53dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1713_l1703_l1697_l1694_l1689_DUPLICATE_53dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1713_l1703_l1697_l1694_l1689_DUPLICATE_53dc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_f825_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_f825_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1707_l1697_l1703_DUPLICATE_f825_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_9eca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_9eca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_9eca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_9eca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1707_l1703_l1697_l1694_l1689_DUPLICATE_9eca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1700_c30_b49e_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1707_c7_c931] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1697_c7_76b8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1701_c22_eddc] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1703_c7_e5bb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;

     -- t8_MUX[uxn_opcodes_h_l1697_c7_76b8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond <= VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond;
     t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue;
     t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output := t8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1707_c7_c931] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_return_output := result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1689_c1_7a1c] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1713_c7_1319] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1707_c7_c931] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_cond;
     tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_return_output := tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1705_c22_3c8e] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1713_c7_1319] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1701_c3_ca3e := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1701_c22_eddc_return_output)),16);
     VAR_result_u16_value_uxn_opcodes_h_l1705_c3_1917 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1705_c22_3c8e_return_output)),16);
     VAR_printf_uxn_opcodes_h_l1690_c3_acb9_uxn_opcodes_h_l1690_c3_acb9_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1689_c1_7a1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1713_c7_1319_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1713_c7_1319_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1707_c7_c931_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1707_c7_c931_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1707_c7_c931_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1701_c3_ca3e;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1705_c3_1917;
     -- result_u16_value_MUX[uxn_opcodes_h_l1703_c7_e5bb] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output := result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1703_c7_e5bb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1697_c7_76b8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;

     -- printf_uxn_opcodes_h_l1690_c3_acb9[uxn_opcodes_h_l1690_c3_acb9] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1690_c3_acb9_uxn_opcodes_h_l1690_c3_acb9_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1690_c3_acb9_uxn_opcodes_h_l1690_c3_acb9_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l1703_c7_e5bb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output := result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1707_c7_c931] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1694_c7_6df0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1703_c7_e5bb] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond;
     tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output := tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1707_c7_c931] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_return_output;

     -- t8_MUX[uxn_opcodes_h_l1694_c7_6df0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond <= VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond;
     t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue;
     t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output := t8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1707_c7_c931_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1707_c7_c931_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1703_c7_e5bb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1697_c7_76b8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output := result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;

     -- t8_MUX[uxn_opcodes_h_l1689_c2_7f74] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond <= VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond;
     t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue;
     t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output := t8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1703_c7_e5bb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1697_c7_76b8] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output := result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1694_c7_6df0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1697_c7_76b8] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_cond;
     tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output := tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1689_c2_7f74] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1697_c7_76b8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1703_c7_e5bb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1694_c7_6df0] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_cond;
     tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output := tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1694_c7_6df0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1697_c7_76b8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1689_c2_7f74] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1694_c7_6df0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1697_c7_76b8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1694_c7_6df0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output := result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1697_c7_76b8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1689_c2_7f74] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1689_c2_7f74] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output := result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1689_c2_7f74] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output := result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1689_c2_7f74] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_cond;
     tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output := tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1694_c7_6df0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1694_c7_6df0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1694_c7_6df0_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1689_c2_7f74] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1689_c2_7f74] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_9969_uxn_opcodes_h_l1685_l1718_DUPLICATE_3ec6 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9969_uxn_opcodes_h_l1685_l1718_DUPLICATE_3ec6_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_9969(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1689_c2_7f74_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9969_uxn_opcodes_h_l1685_l1718_DUPLICATE_3ec6_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9969_uxn_opcodes_h_l1685_l1718_DUPLICATE_3ec6_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
