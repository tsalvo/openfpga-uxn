-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity sta_0CLK_bce25fe8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sta_0CLK_bce25fe8;
architecture arch of sta_0CLK_bce25fe8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2315_c6_9fe4]
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2315_c2_1128]
signal n8_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2315_c2_1128]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c2_1128]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c2_1128]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2315_c2_1128]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c2_1128]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2315_c2_1128]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2315_c2_1128]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2315_c2_1128]
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2315_c2_1128]
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2315_c2_1128]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2315_c2_1128]
signal t16_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2328_c11_abd8]
signal BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2328_c7_e86c]
signal n8_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2328_c7_e86c]
signal result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2328_c7_e86c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2328_c7_e86c]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2328_c7_e86c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2328_c7_e86c]
signal result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2328_c7_e86c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l2328_c7_e86c]
signal t16_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2331_c11_443f]
signal BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2331_c7_7153]
signal n8_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2331_c7_7153]
signal result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2331_c7_7153]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2331_c7_7153]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2331_c7_7153]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2331_c7_7153]
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2331_c7_7153]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l2331_c7_7153]
signal t16_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2333_c3_2dbc]
signal CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2336_c11_eb3f]
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2336_c7_32eb]
signal n8_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2336_c7_32eb]
signal result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2336_c7_32eb]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2336_c7_32eb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2336_c7_32eb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2336_c7_32eb]
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2336_c7_32eb]
signal t16_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2337_c3_4fea]
signal BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2339_c11_45e1]
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2339_c7_8150]
signal n8_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2339_c7_8150]
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2339_c7_8150]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2339_c7_8150]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2339_c7_8150]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2339_c7_8150]
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2341_c30_c2b6]
signal sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_return_output : signed(3 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_42c1( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u16_value := ref_toks_8;
      base.u8_value := ref_toks_9;
      base.is_vram_write := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4
BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_left,
BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_right,
BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output);

-- n8_MUX_uxn_opcodes_h_l2315_c2_1128
n8_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
n8_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
n8_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
n8_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128
result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128
result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128
result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128
result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- t16_MUX_uxn_opcodes_h_l2315_c2_1128
t16_MUX_uxn_opcodes_h_l2315_c2_1128 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2315_c2_1128_cond,
t16_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue,
t16_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse,
t16_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8
BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_left,
BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_right,
BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output);

-- n8_MUX_uxn_opcodes_h_l2328_c7_e86c
n8_MUX_uxn_opcodes_h_l2328_c7_e86c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2328_c7_e86c_cond,
n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue,
n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse,
n8_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c
result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond,
result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c
result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c
result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c
result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output);

-- t16_MUX_uxn_opcodes_h_l2328_c7_e86c
t16_MUX_uxn_opcodes_h_l2328_c7_e86c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2328_c7_e86c_cond,
t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue,
t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse,
t16_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_left,
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_right,
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output);

-- n8_MUX_uxn_opcodes_h_l2331_c7_7153
n8_MUX_uxn_opcodes_h_l2331_c7_7153 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2331_c7_7153_cond,
n8_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue,
n8_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse,
n8_MUX_uxn_opcodes_h_l2331_c7_7153_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153
result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond,
result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153
result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153
result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond,
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_return_output);

-- t16_MUX_uxn_opcodes_h_l2331_c7_7153
t16_MUX_uxn_opcodes_h_l2331_c7_7153 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2331_c7_7153_cond,
t16_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue,
t16_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse,
t16_MUX_uxn_opcodes_h_l2331_c7_7153_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc
CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_x,
CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_left,
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_right,
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output);

-- n8_MUX_uxn_opcodes_h_l2336_c7_32eb
n8_MUX_uxn_opcodes_h_l2336_c7_32eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2336_c7_32eb_cond,
n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue,
n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse,
n8_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb
result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond,
result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb
result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb
result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond,
result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output);

-- t16_MUX_uxn_opcodes_h_l2336_c7_32eb
t16_MUX_uxn_opcodes_h_l2336_c7_32eb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2336_c7_32eb_cond,
t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue,
t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse,
t16_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea
BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_left,
BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_right,
BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_left,
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_right,
BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output);

-- n8_MUX_uxn_opcodes_h_l2339_c7_8150
n8_MUX_uxn_opcodes_h_l2339_c7_8150 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2339_c7_8150_cond,
n8_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue,
n8_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse,
n8_MUX_uxn_opcodes_h_l2339_c7_8150_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150
result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond,
result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150
result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond,
result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6
sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_ins,
sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_x,
sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_y,
sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output,
 n8_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 t16_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output,
 n8_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output,
 t16_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output,
 n8_MUX_uxn_opcodes_h_l2331_c7_7153_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_return_output,
 t16_MUX_uxn_opcodes_h_l2331_c7_7153_return_output,
 CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output,
 n8_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output,
 t16_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output,
 n8_MUX_uxn_opcodes_h_l2339_c7_8150_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output,
 sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2320_c3_e517 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2325_c3_cc02 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2329_c3_4953 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2334_c3_d463 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2331_c7_7153_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_d69e_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_8c09_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0b8e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0bc5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_1e3e_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2337_l2332_DUPLICATE_f2f0_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l2348_l2310_DUPLICATE_4fad_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2325_c3_cc02 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2325_c3_cc02;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2334_c3_d463 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2334_c3_d463;
     VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_right := to_unsigned(3, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_y := resize(to_signed(-3, 3), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_right := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2320_c3_e517 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2320_c3_e517;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2329_c3_4953 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2329_c3_4953;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_left := t16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse := t16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0bc5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0bc5_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2339_c11_45e1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2315_c6_9fe4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2315_c2_1128_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2331_c11_443f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2337_l2332_DUPLICATE_f2f0 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2337_l2332_DUPLICATE_f2f0_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_8c09 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_8c09_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2328_c11_abd8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0b8e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0b8e_return_output := result.is_opc_done;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2331_c7_7153] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2331_c7_7153_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_1e3e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_1e3e_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2336_c11_eb3f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2341_c30_c2b6] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_ins;
     sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_x;
     sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_return_output := sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2315_c2_1128_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_d69e LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_d69e_return_output := result.u16_value;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2315_c2_1128_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2315_c2_1128_return_output := result.is_vram_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c6_9fe4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2328_c11_abd8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_443f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_eb3f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2339_c11_45e1_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2337_l2332_DUPLICATE_f2f0_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2337_l2332_DUPLICATE_f2f0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_1e3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_1e3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_1e3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_1e3e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_d69e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_d69e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_d69e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_d69e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_d69e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0b8e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0b8e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0b8e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0b8e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0bc5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0bc5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0bc5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2331_l2336_l2328_l2339_DUPLICATE_0bc5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_8c09_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_8c09_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_8c09_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_8c09_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2336_l2331_l2328_l2315_l2339_DUPLICATE_8c09_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2315_c2_1128_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2315_c2_1128_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2315_c2_1128_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2315_c2_1128_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2331_c7_7153_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2341_c30_c2b6_return_output;
     -- BIN_OP_OR[uxn_opcodes_h_l2337_c3_4fea] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_left;
     BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_return_output := BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2331_c7_7153] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2339_c7_8150] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2339_c7_8150] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2339_c7_8150] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2333_c3_2dbc] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_return_output := CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2339_c7_8150] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output := result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2339_c7_8150] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output := result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;

     -- n8_MUX[uxn_opcodes_h_l2339_c7_8150] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2339_c7_8150_cond <= VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_cond;
     n8_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_iftrue;
     n8_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_return_output := n8_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2337_c3_4fea_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2333_c3_2dbc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2339_c7_8150_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2336_c7_32eb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2336_c7_32eb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2328_c7_e86c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2336_c7_32eb] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2336_c7_32eb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output := result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;

     -- n8_MUX[uxn_opcodes_h_l2336_c7_32eb] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2336_c7_32eb_cond <= VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_cond;
     n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue;
     n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output := n8_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2336_c7_32eb] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output := result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;

     -- t16_MUX[uxn_opcodes_h_l2336_c7_32eb] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2336_c7_32eb_cond <= VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_cond;
     t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iftrue;
     t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output := t16_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2336_c7_32eb_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2331_c7_7153] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output := result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2331_c7_7153] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2331_c7_7153] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- t16_MUX[uxn_opcodes_h_l2331_c7_7153] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2331_c7_7153_cond <= VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_cond;
     t16_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue;
     t16_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_return_output := t16_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;

     -- n8_MUX[uxn_opcodes_h_l2331_c7_7153] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2331_c7_7153_cond <= VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_cond;
     n8_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue;
     n8_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_return_output := n8_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2331_c7_7153] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2331_c7_7153] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output := result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2331_c7_7153_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2328_c7_e86c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;

     -- t16_MUX[uxn_opcodes_h_l2328_c7_e86c] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2328_c7_e86c_cond <= VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_cond;
     t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue;
     t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output := t16_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2328_c7_e86c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output := result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2328_c7_e86c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2328_c7_e86c] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2328_c7_e86c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2328_c7_e86c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_cond;
     n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue;
     n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output := n8_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2328_c7_e86c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2328_c7_e86c_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- t16_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     t16_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     t16_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := t16_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- n8_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     n8_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     n8_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := n8_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c2_1128] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2315_c2_1128_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l2348_l2310_DUPLICATE_4fad LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l2348_l2310_DUPLICATE_4fad_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_42c1(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c2_1128_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2315_c2_1128_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l2348_l2310_DUPLICATE_4fad_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_42c1_uxn_opcodes_h_l2348_l2310_DUPLICATE_4fad_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
