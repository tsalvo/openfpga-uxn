-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity and_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end and_0CLK_64d180f1;
architecture arch of and_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l921_c6_0934]
signal BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l921_c2_97aa]
signal n8_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l921_c2_97aa]
signal result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l921_c2_97aa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l921_c2_97aa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l921_c2_97aa]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l921_c2_97aa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l921_c2_97aa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l921_c2_97aa]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l921_c2_97aa]
signal result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l921_c2_97aa]
signal result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l921_c2_97aa]
signal t8_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l934_c11_b714]
signal BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l934_c7_448a]
signal n8_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l934_c7_448a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l934_c7_448a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l934_c7_448a]
signal result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l934_c7_448a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l934_c7_448a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l934_c7_448a]
signal t8_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l937_c11_a03e]
signal BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l937_c7_06d8]
signal n8_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l937_c7_06d8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l937_c7_06d8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l937_c7_06d8]
signal result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l937_c7_06d8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l937_c7_06d8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l937_c7_06d8]
signal t8_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l940_c11_4f2a]
signal BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l940_c7_c71e]
signal n8_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l940_c7_c71e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l940_c7_c71e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l940_c7_c71e]
signal result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l940_c7_c71e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l940_c7_c71e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l942_c30_a2c4]
signal sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l945_c21_740a]
signal BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a47b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934
BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_left,
BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_right,
BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output);

-- n8_MUX_uxn_opcodes_h_l921_c2_97aa
n8_MUX_uxn_opcodes_h_l921_c2_97aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l921_c2_97aa_cond,
n8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue,
n8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse,
n8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa
result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa
result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa
result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa
result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa
result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa
result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_cond,
result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa
result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

-- t8_MUX_uxn_opcodes_h_l921_c2_97aa
t8_MUX_uxn_opcodes_h_l921_c2_97aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l921_c2_97aa_cond,
t8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue,
t8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse,
t8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714
BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_left,
BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_right,
BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output);

-- n8_MUX_uxn_opcodes_h_l934_c7_448a
n8_MUX_uxn_opcodes_h_l934_c7_448a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l934_c7_448a_cond,
n8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue,
n8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse,
n8_MUX_uxn_opcodes_h_l934_c7_448a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a
result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a
result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a
result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_cond,
result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a
result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_return_output);

-- t8_MUX_uxn_opcodes_h_l934_c7_448a
t8_MUX_uxn_opcodes_h_l934_c7_448a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l934_c7_448a_cond,
t8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue,
t8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse,
t8_MUX_uxn_opcodes_h_l934_c7_448a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e
BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_left,
BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_right,
BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output);

-- n8_MUX_uxn_opcodes_h_l937_c7_06d8
n8_MUX_uxn_opcodes_h_l937_c7_06d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l937_c7_06d8_cond,
n8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue,
n8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse,
n8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8
result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8
result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8
result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_cond,
result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8
result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_return_output);

-- t8_MUX_uxn_opcodes_h_l937_c7_06d8
t8_MUX_uxn_opcodes_h_l937_c7_06d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l937_c7_06d8_cond,
t8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue,
t8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse,
t8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a
BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_left,
BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_right,
BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output);

-- n8_MUX_uxn_opcodes_h_l940_c7_c71e
n8_MUX_uxn_opcodes_h_l940_c7_c71e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l940_c7_c71e_cond,
n8_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue,
n8_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse,
n8_MUX_uxn_opcodes_h_l940_c7_c71e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e
result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e
result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e
result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_cond,
result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e
result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_return_output);

-- sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4
sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_ins,
sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_x,
sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_y,
sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l945_c21_740a
BIN_OP_AND_uxn_opcodes_h_l945_c21_740a : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_left,
BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_right,
BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output,
 n8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
 t8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output,
 n8_MUX_uxn_opcodes_h_l934_c7_448a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_return_output,
 t8_MUX_uxn_opcodes_h_l934_c7_448a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output,
 n8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_return_output,
 t8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output,
 n8_MUX_uxn_opcodes_h_l940_c7_c71e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_return_output,
 sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_return_output,
 BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l926_c3_beac : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l931_c3_cc19 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l935_c3_9718 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l944_c3_a713 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l934_l937_l940_l921_DUPLICATE_fa6f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_47f0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_d548_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_f5ec_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l937_l940_DUPLICATE_90c4_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l949_l917_DUPLICATE_1c80_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l931_c3_cc19 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l931_c3_cc19;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l935_c3_9718 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l935_c3_9718;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_right := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l926_c3_beac := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l926_c3_beac;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l944_c3_a713 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l944_c3_a713;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l940_c11_4f2a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_left;
     BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output := BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l921_c2_97aa_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l921_c6_0934] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_left;
     BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output := BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_d548 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_d548_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l942_c30_a2c4] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_ins;
     sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_x <= VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_x;
     sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_y <= VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_return_output := sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l945_c21_740a] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_left;
     BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_return_output := BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l921_c2_97aa_return_output := result.is_stack_index_flipped;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l921_c2_97aa_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l937_c11_a03e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_left;
     BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output := BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l934_c11_b714] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_left;
     BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output := BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l934_l937_l940_l921_DUPLICATE_fa6f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l934_l937_l940_l921_DUPLICATE_fa6f_return_output := result.u8_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l937_l940_DUPLICATE_90c4 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l937_l940_DUPLICATE_90c4_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_f5ec LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_f5ec_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l921_c2_97aa_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_47f0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_47f0_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l945_c21_740a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l921_c6_0934_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l934_c11_b714_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l937_c11_a03e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l940_c11_4f2a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_d548_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_d548_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_d548_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_47f0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_47f0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_47f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_f5ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_f5ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l934_l937_l940_DUPLICATE_f5ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l937_l940_DUPLICATE_90c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l937_l940_DUPLICATE_90c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l934_l937_l940_l921_DUPLICATE_fa6f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l934_l937_l940_l921_DUPLICATE_fa6f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l934_l937_l940_l921_DUPLICATE_fa6f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l934_l937_l940_l921_DUPLICATE_fa6f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l921_c2_97aa_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l921_c2_97aa_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l921_c2_97aa_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l921_c2_97aa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l942_c30_a2c4_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l940_c7_c71e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;

     -- t8_MUX[uxn_opcodes_h_l937_c7_06d8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l937_c7_06d8_cond <= VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_cond;
     t8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue;
     t8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output := t8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;

     -- n8_MUX[uxn_opcodes_h_l940_c7_c71e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l940_c7_c71e_cond <= VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_cond;
     n8_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue;
     n8_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_return_output := n8_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l940_c7_c71e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_return_output := result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l940_c7_c71e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l940_c7_c71e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l940_c7_c71e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l940_c7_c71e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;
     -- t8_MUX[uxn_opcodes_h_l934_c7_448a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l934_c7_448a_cond <= VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_cond;
     t8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue;
     t8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_return_output := t8_MUX_uxn_opcodes_h_l934_c7_448a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l937_c7_06d8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l937_c7_06d8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l937_c7_06d8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;

     -- n8_MUX[uxn_opcodes_h_l937_c7_06d8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l937_c7_06d8_cond <= VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_cond;
     n8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue;
     n8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output := n8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l937_c7_06d8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_return_output := result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l937_c7_06d8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l937_c7_06d8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse := VAR_t8_MUX_uxn_opcodes_h_l934_c7_448a_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l934_c7_448a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l934_c7_448a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_return_output;

     -- t8_MUX[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l921_c2_97aa_cond <= VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_cond;
     t8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue;
     t8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output := t8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l934_c7_448a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_return_output := result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_return_output;

     -- n8_MUX[uxn_opcodes_h_l934_c7_448a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l934_c7_448a_cond <= VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_cond;
     n8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_iftrue;
     n8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_return_output := n8_MUX_uxn_opcodes_h_l934_c7_448a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l934_c7_448a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l934_c7_448a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse := VAR_n8_MUX_uxn_opcodes_h_l934_c7_448a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l934_c7_448a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l934_c7_448a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l934_c7_448a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l934_c7_448a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l934_c7_448a_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;
     -- n8_MUX[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l921_c2_97aa_cond <= VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_cond;
     n8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue;
     n8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output := n8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_return_output := result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l921_c2_97aa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l921_c2_97aa_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l949_l917_DUPLICATE_1c80 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l949_l917_DUPLICATE_1c80_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a47b(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l921_c2_97aa_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l921_c2_97aa_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l949_l917_DUPLICATE_1c80_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l949_l917_DUPLICATE_1c80_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
