-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity gth_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_226c8821;
architecture arch of gth_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1826_c6_2dd9]
signal BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1826_c2_787d]
signal t8_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1826_c2_787d]
signal n8_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1826_c2_787d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1826_c2_787d]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1826_c2_787d]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1826_c2_787d]
signal result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1826_c2_787d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1826_c2_787d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1826_c2_787d]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1826_c2_787d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1826_c2_787d]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1839_c11_a68a]
signal BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1839_c7_db5e]
signal t8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1839_c7_db5e]
signal n8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1839_c7_db5e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1839_c7_db5e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1839_c7_db5e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1839_c7_db5e]
signal result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1839_c7_db5e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1842_c11_d6c7]
signal BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1842_c7_42f9]
signal t8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1842_c7_42f9]
signal n8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1842_c7_42f9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1842_c7_42f9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1842_c7_42f9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1842_c7_42f9]
signal result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1842_c7_42f9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1845_c11_4e1f]
signal BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1845_c7_b38c]
signal n8_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1845_c7_b38c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1845_c7_b38c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1845_c7_b38c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1845_c7_b38c]
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1845_c7_b38c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1847_c30_f9de]
signal sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1850_c21_bf4e]
signal BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1850_c21_3c37]
signal MUX_uxn_opcodes_h_l1850_c21_3c37_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1850_c21_3c37_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1850_c21_3c37_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1850_c21_3c37_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_188e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_ram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9
BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_left,
BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_right,
BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output);

-- t8_MUX_uxn_opcodes_h_l1826_c2_787d
t8_MUX_uxn_opcodes_h_l1826_c2_787d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1826_c2_787d_cond,
t8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue,
t8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse,
t8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

-- n8_MUX_uxn_opcodes_h_l1826_c2_787d
n8_MUX_uxn_opcodes_h_l1826_c2_787d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1826_c2_787d_cond,
n8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue,
n8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse,
n8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d
result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d
result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d
result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d
result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a
BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_left,
BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_right,
BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output);

-- t8_MUX_uxn_opcodes_h_l1839_c7_db5e
t8_MUX_uxn_opcodes_h_l1839_c7_db5e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond,
t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue,
t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse,
t8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output);

-- n8_MUX_uxn_opcodes_h_l1839_c7_db5e
n8_MUX_uxn_opcodes_h_l1839_c7_db5e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond,
n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue,
n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse,
n8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e
result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e
result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e
result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7
BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_left,
BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_right,
BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output);

-- t8_MUX_uxn_opcodes_h_l1842_c7_42f9
t8_MUX_uxn_opcodes_h_l1842_c7_42f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond,
t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue,
t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse,
t8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output);

-- n8_MUX_uxn_opcodes_h_l1842_c7_42f9
n8_MUX_uxn_opcodes_h_l1842_c7_42f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond,
n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue,
n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse,
n8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9
result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9
result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9
result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_left,
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_right,
BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output);

-- n8_MUX_uxn_opcodes_h_l1845_c7_b38c
n8_MUX_uxn_opcodes_h_l1845_c7_b38c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1845_c7_b38c_cond,
n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue,
n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse,
n8_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de
sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_ins,
sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_x,
sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_y,
sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e
BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_left,
BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_right,
BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_return_output);

-- MUX_uxn_opcodes_h_l1850_c21_3c37
MUX_uxn_opcodes_h_l1850_c21_3c37 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1850_c21_3c37_cond,
MUX_uxn_opcodes_h_l1850_c21_3c37_iftrue,
MUX_uxn_opcodes_h_l1850_c21_3c37_iffalse,
MUX_uxn_opcodes_h_l1850_c21_3c37_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output,
 t8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
 n8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output,
 t8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output,
 n8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output,
 t8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output,
 n8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output,
 n8_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output,
 sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_return_output,
 MUX_uxn_opcodes_h_l1850_c21_3c37_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1831_c3_99b5 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1836_c3_1833 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1840_c3_b4b0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1849_c3_09c9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1842_l1826_l1845_l1839_DUPLICATE_b5f0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_99ec_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_8f53_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_1b59_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1842_l1845_DUPLICATE_2e73_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1854_l1822_DUPLICATE_6378_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_right := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1849_c3_09c9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1849_c3_09c9;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1836_c3_1833 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1836_c3_1833;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1840_c3_b4b0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1840_c3_b4b0;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_y := resize(to_signed(-1, 2), 4);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1831_c3_99b5 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1831_c3_99b5;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse := t8;
     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1826_c2_787d_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_1b59 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_1b59_return_output := result.is_opc_done;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1826_c2_787d_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1842_l1826_l1845_l1839_DUPLICATE_b5f0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1842_l1826_l1845_l1839_DUPLICATE_b5f0_return_output := result.u8_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1842_l1845_DUPLICATE_2e73 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1842_l1845_DUPLICATE_2e73_return_output := result.stack_address_sp_offset;

     -- BIN_OP_GT[uxn_opcodes_h_l1850_c21_bf4e] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_left;
     BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_return_output := BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1845_c11_4e1f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1826_c2_787d_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1826_c6_2dd9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1839_c11_a68a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1826_c2_787d_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l1847_c30_f9de] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_ins;
     sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_x;
     sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_return_output := sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_99ec LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_99ec_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_8f53 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_8f53_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1842_c11_d6c7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1826_c6_2dd9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1839_c11_a68a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1842_c11_d6c7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1845_c11_4e1f_return_output;
     VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1850_c21_bf4e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_99ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_99ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_99ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_1b59_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_1b59_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_1b59_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_8f53_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_8f53_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1842_l1845_l1839_DUPLICATE_8f53_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1842_l1845_DUPLICATE_2e73_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1842_l1845_DUPLICATE_2e73_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1842_l1826_l1845_l1839_DUPLICATE_b5f0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1842_l1826_l1845_l1839_DUPLICATE_b5f0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1842_l1826_l1845_l1839_DUPLICATE_b5f0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1842_l1826_l1845_l1839_DUPLICATE_b5f0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1826_c2_787d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1826_c2_787d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1826_c2_787d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1826_c2_787d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1847_c30_f9de_return_output;
     -- n8_MUX[uxn_opcodes_h_l1845_c7_b38c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1845_c7_b38c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_cond;
     n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue;
     n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output := n8_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;

     -- t8_MUX[uxn_opcodes_h_l1842_c7_42f9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond <= VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond;
     t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue;
     t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output := t8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1845_c7_b38c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1845_c7_b38c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1845_c7_b38c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1845_c7_b38c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;

     -- MUX[uxn_opcodes_h_l1850_c21_3c37] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1850_c21_3c37_cond <= VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_cond;
     MUX_uxn_opcodes_h_l1850_c21_3c37_iftrue <= VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_iftrue;
     MUX_uxn_opcodes_h_l1850_c21_3c37_iffalse <= VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_return_output := MUX_uxn_opcodes_h_l1850_c21_3c37_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue := VAR_MUX_uxn_opcodes_h_l1850_c21_3c37_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1842_c7_42f9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1842_c7_42f9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1845_c7_b38c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1839_c7_db5e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond;
     t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue;
     t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output := t8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;

     -- n8_MUX[uxn_opcodes_h_l1842_c7_42f9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond <= VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_cond;
     n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue;
     n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output := n8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1842_c7_42f9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1842_c7_42f9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1845_c7_b38c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1839_c7_db5e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1839_c7_db5e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1839_c7_db5e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1842_c7_42f9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;

     -- t8_MUX[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1826_c2_787d_cond <= VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_cond;
     t8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue;
     t8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output := t8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;

     -- n8_MUX[uxn_opcodes_h_l1839_c7_db5e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond <= VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_cond;
     n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue;
     n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output := n8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1839_c7_db5e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1842_c7_42f9_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;

     -- n8_MUX[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1826_c2_787d_cond <= VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_cond;
     n8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue;
     n8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output := n8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1839_c7_db5e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1839_c7_db5e_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1826_c2_787d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1854_l1822_DUPLICATE_6378 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1854_l1822_DUPLICATE_6378_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_188e(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1826_c2_787d_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1826_c2_787d_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1854_l1822_DUPLICATE_6378_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1854_l1822_DUPLICATE_6378_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
