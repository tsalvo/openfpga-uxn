-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity lth_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_85d5529e;
architecture arch of lth_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1800_c6_cd0e]
signal BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1800_c1_aba9]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1800_c2_3869]
signal t8_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1800_c2_3869]
signal n8_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1800_c2_3869]
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1800_c2_3869]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1800_c2_3869]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1800_c2_3869]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1800_c2_3869]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1800_c2_3869]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l1801_c3_d38e[uxn_opcodes_h_l1801_c3_d38e]
signal printf_uxn_opcodes_h_l1801_c3_d38e_uxn_opcodes_h_l1801_c3_d38e_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1805_c11_303c]
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1805_c7_8eba]
signal t8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1805_c7_8eba]
signal n8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1805_c7_8eba]
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1805_c7_8eba]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1805_c7_8eba]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1805_c7_8eba]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1805_c7_8eba]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1805_c7_8eba]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1808_c11_828b]
signal BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1808_c7_1cfb]
signal t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1808_c7_1cfb]
signal n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1808_c7_1cfb]
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1808_c7_1cfb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1808_c7_1cfb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1808_c7_1cfb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1808_c7_1cfb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1808_c7_1cfb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1811_c11_c2d7]
signal BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1811_c7_7654]
signal n8_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1811_c7_7654]
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1811_c7_7654]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1811_c7_7654]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1811_c7_7654]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1811_c7_7654]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1811_c7_7654]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1814_c30_11b2]
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l1817_c21_8b2d]
signal BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1817_c21_dfde]
signal MUX_uxn_opcodes_h_l1817_c21_dfde_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1817_c21_dfde_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1817_c21_dfde_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1817_c21_dfde_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1819_c11_ba6f]
signal BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1819_c7_5885]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1819_c7_5885]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1819_c7_5885]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_left,
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_right,
BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_return_output);

-- t8_MUX_uxn_opcodes_h_l1800_c2_3869
t8_MUX_uxn_opcodes_h_l1800_c2_3869 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1800_c2_3869_cond,
t8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue,
t8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse,
t8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output);

-- n8_MUX_uxn_opcodes_h_l1800_c2_3869
n8_MUX_uxn_opcodes_h_l1800_c2_3869 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1800_c2_3869_cond,
n8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue,
n8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse,
n8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_cond,
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output);

-- printf_uxn_opcodes_h_l1801_c3_d38e_uxn_opcodes_h_l1801_c3_d38e
printf_uxn_opcodes_h_l1801_c3_d38e_uxn_opcodes_h_l1801_c3_d38e : entity work.printf_uxn_opcodes_h_l1801_c3_d38e_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1801_c3_d38e_uxn_opcodes_h_l1801_c3_d38e_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_left,
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_right,
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output);

-- t8_MUX_uxn_opcodes_h_l1805_c7_8eba
t8_MUX_uxn_opcodes_h_l1805_c7_8eba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond,
t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue,
t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse,
t8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output);

-- n8_MUX_uxn_opcodes_h_l1805_c7_8eba
n8_MUX_uxn_opcodes_h_l1805_c7_8eba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond,
n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue,
n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse,
n8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_cond,
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_left,
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_right,
BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output);

-- t8_MUX_uxn_opcodes_h_l1808_c7_1cfb
t8_MUX_uxn_opcodes_h_l1808_c7_1cfb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond,
t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue,
t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse,
t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output);

-- n8_MUX_uxn_opcodes_h_l1808_c7_1cfb
n8_MUX_uxn_opcodes_h_l1808_c7_1cfb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond,
n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue,
n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse,
n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond,
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_left,
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_right,
BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output);

-- n8_MUX_uxn_opcodes_h_l1811_c7_7654
n8_MUX_uxn_opcodes_h_l1811_c7_7654 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1811_c7_7654_cond,
n8_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue,
n8_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse,
n8_MUX_uxn_opcodes_h_l1811_c7_7654_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_cond,
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2
sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_ins,
sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_x,
sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_y,
sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d
BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_left,
BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_right,
BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_return_output);

-- MUX_uxn_opcodes_h_l1817_c21_dfde
MUX_uxn_opcodes_h_l1817_c21_dfde : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1817_c21_dfde_cond,
MUX_uxn_opcodes_h_l1817_c21_dfde_iftrue,
MUX_uxn_opcodes_h_l1817_c21_dfde_iffalse,
MUX_uxn_opcodes_h_l1817_c21_dfde_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_left,
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_right,
BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_return_output,
 t8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
 n8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output,
 t8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output,
 n8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output,
 t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output,
 n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output,
 n8_MUX_uxn_opcodes_h_l1811_c7_7654_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output,
 sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_return_output,
 BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_return_output,
 MUX_uxn_opcodes_h_l1817_c21_dfde_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_8978 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1801_c3_d38e_uxn_opcodes_h_l1801_c3_d38e_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1806_c3_9c1f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1816_c3_71e5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_7287_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_6e9b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_fee5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_1549_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1811_DUPLICATE_60ef_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1808_l1811_DUPLICATE_28de_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1796_l1825_DUPLICATE_5273_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1816_c3_71e5 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1816_c3_71e5;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_8978 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_8978;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1806_c3_9c1f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1806_c3_9c1f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_right := to_unsigned(4, 3);
     VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1811_c11_c2d7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_7287 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_7287_return_output := result.u8_value;

     -- BIN_OP_LT[uxn_opcodes_h_l1817_c21_8b2d] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_left;
     BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_return_output := BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_fee5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_fee5_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1800_c6_cd0e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_6e9b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_6e9b_return_output := result.is_sp_shift;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_1549 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_1549_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1805_c11_303c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1814_c30_11b2] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_ins;
     sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_x;
     sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_return_output := sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1819_c11_ba6f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1808_l1811_DUPLICATE_28de LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1808_l1811_DUPLICATE_28de_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1808_c11_828b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1811_DUPLICATE_60ef LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1811_DUPLICATE_60ef_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1800_c6_cd0e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_303c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1808_c11_828b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1811_c11_c2d7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1819_c11_ba6f_return_output;
     VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l1817_c21_8b2d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_1549_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_1549_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_1549_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_1549_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1811_DUPLICATE_60ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1811_DUPLICATE_60ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1811_DUPLICATE_60ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1811_DUPLICATE_60ef_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_6e9b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_6e9b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_6e9b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_6e9b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_fee5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_fee5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_fee5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1805_l1819_l1808_l1800_DUPLICATE_fee5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1808_l1811_DUPLICATE_28de_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1808_l1811_DUPLICATE_28de_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_7287_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_7287_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_7287_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1805_l1808_l1800_l1811_DUPLICATE_7287_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1814_c30_11b2_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1811_c7_7654] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;

     -- t8_MUX[uxn_opcodes_h_l1808_c7_1cfb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond <= VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond;
     t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue;
     t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output := t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1800_c1_aba9] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_return_output;

     -- n8_MUX[uxn_opcodes_h_l1811_c7_7654] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1811_c7_7654_cond <= VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_cond;
     n8_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue;
     n8_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_return_output := n8_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1819_c7_5885] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1819_c7_5885] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1811_c7_7654] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;

     -- MUX[uxn_opcodes_h_l1817_c21_dfde] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1817_c21_dfde_cond <= VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_cond;
     MUX_uxn_opcodes_h_l1817_c21_dfde_iftrue <= VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_iftrue;
     MUX_uxn_opcodes_h_l1817_c21_dfde_iffalse <= VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_return_output := MUX_uxn_opcodes_h_l1817_c21_dfde_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1819_c7_5885] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue := VAR_MUX_uxn_opcodes_h_l1817_c21_dfde_return_output;
     VAR_printf_uxn_opcodes_h_l1801_c3_d38e_uxn_opcodes_h_l1801_c3_d38e_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1800_c1_aba9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1819_c7_5885_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1819_c7_5885_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1819_c7_5885_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1808_c7_1cfb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1808_c7_1cfb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1811_c7_7654] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1811_c7_7654] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1811_c7_7654] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_return_output := result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;

     -- n8_MUX[uxn_opcodes_h_l1808_c7_1cfb] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond <= VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond;
     n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue;
     n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output := n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;

     -- printf_uxn_opcodes_h_l1801_c3_d38e[uxn_opcodes_h_l1801_c3_d38e] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1801_c3_d38e_uxn_opcodes_h_l1801_c3_d38e_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1801_c3_d38e_uxn_opcodes_h_l1801_c3_d38e_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1811_c7_7654] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;

     -- t8_MUX[uxn_opcodes_h_l1805_c7_8eba] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond <= VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond;
     t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue;
     t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output := t8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1811_c7_7654_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1805_c7_8eba] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1805_c7_8eba] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;

     -- n8_MUX[uxn_opcodes_h_l1805_c7_8eba] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond <= VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_cond;
     n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue;
     n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output := n8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;

     -- t8_MUX[uxn_opcodes_h_l1800_c2_3869] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1800_c2_3869_cond <= VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_cond;
     t8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue;
     t8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output := t8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1808_c7_1cfb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1808_c7_1cfb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1808_c7_1cfb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1808_c7_1cfb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output := result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1808_c7_1cfb_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1805_c7_8eba] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1800_c2_3869] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1805_c7_8eba] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output := result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;

     -- n8_MUX[uxn_opcodes_h_l1800_c2_3869] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1800_c2_3869_cond <= VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_cond;
     n8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue;
     n8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output := n8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1800_c2_3869] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1805_c7_8eba] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1805_c7_8eba] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1800_c2_3869_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1805_c7_8eba_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1800_c2_3869] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1800_c2_3869] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1800_c2_3869] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_return_output := result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1800_c2_3869] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1796_l1825_DUPLICATE_5273 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1796_l1825_DUPLICATE_5273_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1800_c2_3869_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1800_c2_3869_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1796_l1825_DUPLICATE_5273_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1796_l1825_DUPLICATE_5273_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
