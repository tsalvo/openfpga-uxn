-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity opc_add_phased_0CLK_c3dfc98c is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_add_phased_0CLK_c3dfc98c;
architecture arch of opc_add_phased_0CLK_c3dfc98c is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l1011_c6_1335]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1011_c1_d713]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1014_c7_547c]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1011_c2_bcdd]
signal t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1011_c2_bcdd]
signal n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1011_c2_bcdd]
signal result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l1012_c12_3ff1]
signal set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1014_c11_b7be]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1014_c1_e729]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1017_c7_7ede]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1014_c7_547c]
signal t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1014_c7_547c]
signal n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1014_c7_547c]
signal result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l1015_c8_555b]
signal t_register_uxn_opcodes_phased_h_l1015_c8_555b_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l1015_c8_555b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1017_c11_3c1a]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1017_c1_9a7f]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1020_c7_eb13]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1017_c7_7ede]
signal t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1017_c7_7ede]
signal n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1017_c7_7ede]
signal result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l1018_c8_ef23]
signal n_register_uxn_opcodes_phased_h_l1018_c8_ef23_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l1018_c8_ef23_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1020_c11_322c]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1020_c1_69a8]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1023_c7_fcde]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1020_c7_eb13]
signal n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1020_c7_eb13]
signal result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l1021_c8_f1f3]
signal n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1023_c11_8795]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1023_c1_cb96]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1026_c7_acd7]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1023_c7_fcde]
signal result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l1024_c3_f338]
signal set_uxn_opcodes_phased_h_l1024_c3_f338_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l1024_c3_f338_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1024_c3_f338_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l1024_c3_f338_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1024_c3_f338_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1024_c3_f338_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1024_c3_f338_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1026_c11_e820]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1026_c1_f6ff]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1026_c7_acd7]
signal result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_phased_h_l1027_c33_cefe]
signal BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_right : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_return_output : unsigned(8 downto 0);

-- put_stack[uxn_opcodes_phased_h_l1027_c3_dc17]
signal put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1029_c11_1722]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1029_c7_8af7]
signal result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335
BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd
t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond,
t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd
n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond,
n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd
result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond,
result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue,
result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse,
result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1
set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1 : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_sp,
set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_k,
set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_mul,
set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_add,
set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be
BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c
t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond,
t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c
n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond,
n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1014_c7_547c
result_MUX_uxn_opcodes_phased_h_l1014_c7_547c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond,
result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue,
result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse,
result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output);

-- t_register_uxn_opcodes_phased_h_l1015_c8_555b
t_register_uxn_opcodes_phased_h_l1015_c8_555b : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l1015_c8_555b_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_index,
t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_ptr,
t_register_uxn_opcodes_phased_h_l1015_c8_555b_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a
BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede
t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond,
t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede
n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond,
n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede
result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond,
result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue,
result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse,
result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output);

-- n_register_uxn_opcodes_phased_h_l1018_c8_ef23
n_register_uxn_opcodes_phased_h_l1018_c8_ef23 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l1018_c8_ef23_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_index,
n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_ptr,
n_register_uxn_opcodes_phased_h_l1018_c8_ef23_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c
BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13
n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond,
n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13
result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond,
result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue,
result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse,
result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output);

-- n_register_uxn_opcodes_phased_h_l1021_c8_f1f3
n_register_uxn_opcodes_phased_h_l1021_c8_f1f3 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_index,
n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_ptr,
n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795
BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde
result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond,
result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue,
result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse,
result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output);

-- set_uxn_opcodes_phased_h_l1024_c3_f338
set_uxn_opcodes_phased_h_l1024_c3_f338 : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l1024_c3_f338_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l1024_c3_f338_sp,
set_uxn_opcodes_phased_h_l1024_c3_f338_stack_index,
set_uxn_opcodes_phased_h_l1024_c3_f338_ins,
set_uxn_opcodes_phased_h_l1024_c3_f338_k,
set_uxn_opcodes_phased_h_l1024_c3_f338_mul,
set_uxn_opcodes_phased_h_l1024_c3_f338_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820
BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7
result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond,
result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue,
result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse,
result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output);

-- BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe
BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe : entity work.BIN_OP_PLUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_left,
BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_right,
BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_return_output);

-- put_stack_uxn_opcodes_phased_h_l1027_c3_dc17
put_stack_uxn_opcodes_phased_h_l1027_c3_dc17 : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_sp,
put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_stack_index,
put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_offset,
put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722
BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7
result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_cond,
result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iftrue,
result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iffalse,
result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 n8,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output,
 result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output,
 set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output,
 result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output,
 t_register_uxn_opcodes_phased_h_l1015_c8_555b_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output,
 result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output,
 n_register_uxn_opcodes_phased_h_l1018_c8_ef23_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output,
 result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output,
 n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output,
 result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_return_output,
 result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output,
 BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_return_output,
 result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_value : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_return_output : unsigned(8 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_right := to_unsigned(2, 2);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_right := to_unsigned(4, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue := to_unsigned(0, 1);
     VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_offset := resize(to_unsigned(0, 1), 8);
     VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_mul := resize(to_unsigned(2, 2), 8);
     VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iffalse := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_mul := resize(to_unsigned(2, 2), 8);
     VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_add := resize(to_signed(-1, 2), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_add := resize(to_signed(-1, 2), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_k := VAR_k;
     VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_left := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iffalse := result;
     VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_ptr := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_index := VAR_stack_index;
     VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_index := VAR_stack_index;
     VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_right := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1014_c11_b7be] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1029_c11_1722] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1017_c11_3c1a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1011_c6_1335] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1026_c11_e820] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1020_c11_322c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_phased_h_l1027_c33_cefe] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_left <= VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_left;
     BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_right <= VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_return_output := BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1023_c11_8795] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1011_c6_1335_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1014_c11_b7be_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1017_c11_3c1a_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1020_c11_322c_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1023_c11_8795_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1026_c11_e820_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1029_c11_1722_return_output;
     VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_value := resize(VAR_BIN_OP_PLUS_uxn_opcodes_phased_h_l1027_c33_cefe_return_output, 8);
     -- result_MUX[uxn_opcodes_phased_h_l1029_c7_8af7] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_cond;
     result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_return_output := result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1014_c7_547c] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1011_c1_d713] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1011_c1_d713_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1029_c7_8af7_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1017_c7_7ede] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output;

     -- set_will_fail[uxn_opcodes_phased_h_l1012_c12_3ff1] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_sp;
     set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_k;
     set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_mul;
     set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_return_output := set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1014_c1_e729] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1026_c7_acd7] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond;
     result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output := result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1014_c1_e729_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l1012_c12_3ff1_return_output;
     -- t_register[uxn_opcodes_phased_h_l1015_c8_555b] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l1015_c8_555b_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_index;
     t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_return_output := t_register_uxn_opcodes_phased_h_l1015_c8_555b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1017_c1_9a7f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1023_c7_fcde] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond;
     result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output := result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1020_c7_eb13] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1017_c1_9a7f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue := VAR_t_register_uxn_opcodes_phased_h_l1015_c8_555b_return_output;
     -- n_register[uxn_opcodes_phased_h_l1018_c8_ef23] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l1018_c8_ef23_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_index;
     n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_return_output := n_register_uxn_opcodes_phased_h_l1018_c8_ef23_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1020_c1_69a8] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1020_c7_eb13] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond;
     result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output := result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1023_c7_fcde] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c7_fcde_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1020_c1_69a8_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue := VAR_n_register_uxn_opcodes_phased_h_l1018_c8_ef23_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output;
     -- t8_MUX[uxn_opcodes_phased_h_l1017_c7_7ede] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond;
     t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output := t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1023_c1_cb96] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_return_output;

     -- n_register[uxn_opcodes_phased_h_l1021_c8_f1f3] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_index;
     n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_return_output := n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1026_c7_acd7] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1017_c7_7ede] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond;
     result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output := result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output;

     -- Submodule level 6
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c7_acd7_return_output;
     VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1023_c1_cb96_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue := VAR_n_register_uxn_opcodes_phased_h_l1021_c8_f1f3_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output;
     -- t8_MUX[uxn_opcodes_phased_h_l1014_c7_547c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond;
     t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output := t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1014_c7_547c] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond;
     result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output := result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1026_c1_f6ff] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l1020_c7_eb13] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_cond;
     n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output := n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output;

     -- set[uxn_opcodes_phased_h_l1024_c3_f338] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l1024_c3_f338_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l1024_c3_f338_sp <= VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_sp;
     set_uxn_opcodes_phased_h_l1024_c3_f338_stack_index <= VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_stack_index;
     set_uxn_opcodes_phased_h_l1024_c3_f338_ins <= VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_ins;
     set_uxn_opcodes_phased_h_l1024_c3_f338_k <= VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_k;
     set_uxn_opcodes_phased_h_l1024_c3_f338_mul <= VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_mul;
     set_uxn_opcodes_phased_h_l1024_c3_f338_add <= VAR_set_uxn_opcodes_phased_h_l1024_c3_f338_add;
     -- Outputs

     -- Submodule level 7
     VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1026_c1_f6ff_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1020_c7_eb13_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1017_c7_7ede] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_cond;
     n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output := n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l1011_c2_bcdd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond;
     t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output := t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1011_c2_bcdd] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond;
     result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output := result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output;

     -- put_stack[uxn_opcodes_phased_h_l1027_c3_dc17] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_sp <= VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_sp;
     put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_stack_index;
     put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_offset <= VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_offset;
     put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_value <= VAR_put_stack_uxn_opcodes_phased_h_l1027_c3_dc17_value;
     -- Outputs

     -- Submodule level 8
     VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1017_c7_7ede_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1014_c7_547c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_cond;
     n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output := n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output;

     -- Submodule level 9
     VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1014_c7_547c_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1011_c2_bcdd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_cond;
     n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output := n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output;

     -- Submodule level 10
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_phased_h_l1011_c2_bcdd_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
