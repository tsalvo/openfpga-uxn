-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 56
entity swp_0CLK_bf6dd460 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end swp_0CLK_bf6dd460;
architecture arch of swp_0CLK_bf6dd460 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2710_c6_2ddf]
signal BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2710_c1_998f]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2710_c2_e9e3]
signal n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2710_c2_e9e3]
signal t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2710_c2_e9e3]
signal result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2710_c2_e9e3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2710_c2_e9e3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2710_c2_e9e3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2710_c2_e9e3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2710_c2_e9e3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(3 downto 0);

-- printf_uxn_opcodes_h_l2711_c3_5029[uxn_opcodes_h_l2711_c3_5029]
signal printf_uxn_opcodes_h_l2711_c3_5029_uxn_opcodes_h_l2711_c3_5029_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2715_c11_bfea]
signal BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2715_c7_2956]
signal n8_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2715_c7_2956]
signal t8_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2715_c7_2956]
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2715_c7_2956]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2715_c7_2956]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2715_c7_2956]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2715_c7_2956]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2715_c7_2956]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2718_c11_de2e]
signal BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2718_c7_98d3]
signal n8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2718_c7_98d3]
signal t8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2718_c7_98d3]
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2718_c7_98d3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2718_c7_98d3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2718_c7_98d3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2718_c7_98d3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2718_c7_98d3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2722_c11_403f]
signal BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2722_c7_1091]
signal n8_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2722_c7_1091]
signal result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2722_c7_1091]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2722_c7_1091]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2722_c7_1091]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2722_c7_1091]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2722_c7_1091]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2725_c11_9576]
signal BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2725_c7_9387]
signal n8_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2725_c7_9387]
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2725_c7_9387]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2725_c7_9387]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2725_c7_9387]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2725_c7_9387]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2725_c7_9387]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2728_c30_6f87]
signal sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2733_c11_b673]
signal BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2733_c7_8f02]
signal result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2733_c7_8f02]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2733_c7_8f02]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2733_c7_8f02]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2733_c7_8f02]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2738_c11_4610]
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2738_c7_f3d0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2738_c7_f3d0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_25e8( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf
BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_left,
BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_right,
BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_return_output);

-- n8_MUX_uxn_opcodes_h_l2710_c2_e9e3
n8_MUX_uxn_opcodes_h_l2710_c2_e9e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond,
n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue,
n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse,
n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output);

-- t8_MUX_uxn_opcodes_h_l2710_c2_e9e3
t8_MUX_uxn_opcodes_h_l2710_c2_e9e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond,
t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue,
t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse,
t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3
result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3
result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3
result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3
result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output);

-- printf_uxn_opcodes_h_l2711_c3_5029_uxn_opcodes_h_l2711_c3_5029
printf_uxn_opcodes_h_l2711_c3_5029_uxn_opcodes_h_l2711_c3_5029 : entity work.printf_uxn_opcodes_h_l2711_c3_5029_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2711_c3_5029_uxn_opcodes_h_l2711_c3_5029_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea
BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_left,
BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_right,
BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output);

-- n8_MUX_uxn_opcodes_h_l2715_c7_2956
n8_MUX_uxn_opcodes_h_l2715_c7_2956 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2715_c7_2956_cond,
n8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue,
n8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse,
n8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output);

-- t8_MUX_uxn_opcodes_h_l2715_c7_2956
t8_MUX_uxn_opcodes_h_l2715_c7_2956 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2715_c7_2956_cond,
t8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue,
t8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse,
t8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956
result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_cond,
result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_left,
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_right,
BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output);

-- n8_MUX_uxn_opcodes_h_l2718_c7_98d3
n8_MUX_uxn_opcodes_h_l2718_c7_98d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond,
n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue,
n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse,
n8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output);

-- t8_MUX_uxn_opcodes_h_l2718_c7_98d3
t8_MUX_uxn_opcodes_h_l2718_c7_98d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond,
t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue,
t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse,
t8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f
BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_left,
BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_right,
BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output);

-- n8_MUX_uxn_opcodes_h_l2722_c7_1091
n8_MUX_uxn_opcodes_h_l2722_c7_1091 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2722_c7_1091_cond,
n8_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue,
n8_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse,
n8_MUX_uxn_opcodes_h_l2722_c7_1091_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091
result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_cond,
result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091
result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091
result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091
result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091
result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_left,
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_right,
BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output);

-- n8_MUX_uxn_opcodes_h_l2725_c7_9387
n8_MUX_uxn_opcodes_h_l2725_c7_9387 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2725_c7_9387_cond,
n8_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue,
n8_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse,
n8_MUX_uxn_opcodes_h_l2725_c7_9387_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_cond,
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87
sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_ins,
sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_x,
sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_y,
sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673
BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_left,
BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_right,
BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02
result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_cond,
result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02
result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02
result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02
result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_left,
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_right,
BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_return_output,
 n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
 t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output,
 n8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output,
 t8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output,
 n8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output,
 t8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output,
 n8_MUX_uxn_opcodes_h_l2722_c7_1091_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output,
 n8_MUX_uxn_opcodes_h_l2725_c7_9387_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_return_output,
 sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2712_c3_b772 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2711_c3_5029_uxn_opcodes_h_l2711_c3_5029_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2716_c3_4ea6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2720_c3_442a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2723_c3_a87e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2730_c3_e551 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2735_c3_a15d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2733_c7_8f02_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_b7a7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2725_DUPLICATE_5ebe_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2738_l2733_DUPLICATE_a5a0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_cd57_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2738_l2733_l2725_DUPLICATE_e94b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2743_l2706_DUPLICATE_25a6_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2720_c3_442a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2720_c3_442a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2735_c3_a15d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2735_c3_a15d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2723_c3_a87e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2723_c3_a87e;
     VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2712_c3_b772 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2712_c3_b772;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2730_c3_e551 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2730_c3_e551;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2716_c3_4ea6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2716_c3_4ea6;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l2728_c30_6f87] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_ins;
     sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_x;
     sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_return_output := sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_cd57 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_cd57_return_output := result.is_sp_shift;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2725_DUPLICATE_5ebe LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2725_DUPLICATE_5ebe_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2722_c11_403f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2738_l2733_l2725_DUPLICATE_e94b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2738_l2733_l2725_DUPLICATE_e94b_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2718_c11_de2e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2733_c7_8f02] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2733_c7_8f02_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2710_c6_2ddf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_left;
     BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output := BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2715_c11_bfea] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_left;
     BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output := BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_b7a7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_b7a7_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2738_c11_4610] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_left;
     BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_return_output := BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2738_l2733_DUPLICATE_a5a0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2738_l2733_DUPLICATE_a5a0_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2733_c11_b673] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_left;
     BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_return_output := BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2725_c11_9576] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_left;
     BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output := BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2710_c6_2ddf_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2715_c11_bfea_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2718_c11_de2e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2722_c11_403f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2725_c11_9576_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2733_c11_b673_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2738_c11_4610_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2725_DUPLICATE_5ebe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2725_DUPLICATE_5ebe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2725_DUPLICATE_5ebe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2725_DUPLICATE_5ebe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2725_DUPLICATE_5ebe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2738_l2733_l2725_DUPLICATE_e94b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2738_l2733_l2725_DUPLICATE_e94b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2738_l2733_l2725_DUPLICATE_e94b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2738_l2733_l2725_DUPLICATE_e94b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2738_l2733_l2725_DUPLICATE_e94b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2738_l2733_l2725_DUPLICATE_e94b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_cd57_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_cd57_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_cd57_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_cd57_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_cd57_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2738_l2733_DUPLICATE_a5a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2738_l2733_DUPLICATE_a5a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2738_l2733_DUPLICATE_a5a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2738_l2733_DUPLICATE_a5a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2738_l2733_DUPLICATE_a5a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2738_l2733_DUPLICATE_a5a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_b7a7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_b7a7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_b7a7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_b7a7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2722_l2718_l2715_l2710_l2733_DUPLICATE_b7a7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2733_c7_8f02_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2728_c30_6f87_return_output;
     -- n8_MUX[uxn_opcodes_h_l2725_c7_9387] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2725_c7_9387_cond <= VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_cond;
     n8_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue;
     n8_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_return_output := n8_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2733_c7_8f02] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2725_c7_9387] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2738_c7_f3d0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output;

     -- t8_MUX[uxn_opcodes_h_l2718_c7_98d3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond <= VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond;
     t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue;
     t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output := t8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2733_c7_8f02] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output := result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2738_c7_f3d0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2733_c7_8f02] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2710_c1_998f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2711_c3_5029_uxn_opcodes_h_l2711_c3_5029_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2710_c1_998f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2738_c7_f3d0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2722_c7_1091] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;

     -- t8_MUX[uxn_opcodes_h_l2715_c7_2956] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2715_c7_2956_cond <= VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_cond;
     t8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue;
     t8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output := t8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2725_c7_9387] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;

     -- n8_MUX[uxn_opcodes_h_l2722_c7_1091] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2722_c7_1091_cond <= VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_cond;
     n8_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue;
     n8_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_return_output := n8_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2725_c7_9387] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_return_output := result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;

     -- printf_uxn_opcodes_h_l2711_c3_5029[uxn_opcodes_h_l2711_c3_5029] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2711_c3_5029_uxn_opcodes_h_l2711_c3_5029_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2711_c3_5029_uxn_opcodes_h_l2711_c3_5029_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2733_c7_8f02] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2725_c7_9387] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2733_c7_8f02] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2733_c7_8f02_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;
     -- t8_MUX[uxn_opcodes_h_l2710_c2_e9e3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond <= VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond;
     t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue;
     t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output := t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2722_c7_1091] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_return_output := result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;

     -- n8_MUX[uxn_opcodes_h_l2718_c7_98d3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond <= VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_cond;
     n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue;
     n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output := n8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2725_c7_9387] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2718_c7_98d3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2725_c7_9387] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2722_c7_1091] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2722_c7_1091] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2725_c7_9387_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2722_c7_1091] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2715_c7_2956] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;

     -- n8_MUX[uxn_opcodes_h_l2715_c7_2956] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2715_c7_2956_cond <= VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_cond;
     n8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue;
     n8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output := n8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2718_c7_98d3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2722_c7_1091] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2718_c7_98d3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2718_c7_98d3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2722_c7_1091_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2710_c2_e9e3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2718_c7_98d3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2718_c7_98d3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2715_c7_2956] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2715_c7_2956] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_return_output := result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;

     -- n8_MUX[uxn_opcodes_h_l2710_c2_e9e3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond <= VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond;
     n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue;
     n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output := n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2715_c7_2956] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2718_c7_98d3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2710_c2_e9e3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2715_c7_2956] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2710_c2_e9e3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2710_c2_e9e3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2715_c7_2956] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2715_c7_2956_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2710_c2_e9e3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2710_c2_e9e3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2743_l2706_DUPLICATE_25a6 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2743_l2706_DUPLICATE_25a6_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_25e8(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2710_c2_e9e3_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2743_l2706_DUPLICATE_25a6_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2743_l2706_DUPLICATE_25a6_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
