-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity neq_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_226c8821;
architecture arch of neq_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1259_c6_8358]
signal BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1259_c2_6935]
signal t8_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1259_c2_6935]
signal n8_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1259_c2_6935]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1259_c2_6935]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1259_c2_6935]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1259_c2_6935]
signal result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1259_c2_6935]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1259_c2_6935]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1259_c2_6935]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1259_c2_6935]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1259_c2_6935]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1272_c11_5503]
signal BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1272_c7_61a7]
signal t8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1272_c7_61a7]
signal n8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1272_c7_61a7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1272_c7_61a7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1272_c7_61a7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1272_c7_61a7]
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1272_c7_61a7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1275_c11_1149]
signal BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1275_c7_bbc3]
signal t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1275_c7_bbc3]
signal n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1275_c7_bbc3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1275_c7_bbc3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1275_c7_bbc3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1275_c7_bbc3]
signal result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1275_c7_bbc3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1278_c11_f038]
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1278_c7_5eb1]
signal n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1278_c7_5eb1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1278_c7_5eb1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1278_c7_5eb1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1278_c7_5eb1]
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1278_c7_5eb1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1280_c30_f0f2]
signal sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1283_c21_69e3]
signal BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1283_c21_7ac7]
signal MUX_uxn_opcodes_h_l1283_c21_7ac7_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1283_c21_7ac7_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1283_c21_7ac7_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1283_c21_7ac7_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_188e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_ram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358
BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_left,
BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_right,
BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output);

-- t8_MUX_uxn_opcodes_h_l1259_c2_6935
t8_MUX_uxn_opcodes_h_l1259_c2_6935 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1259_c2_6935_cond,
t8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue,
t8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse,
t8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

-- n8_MUX_uxn_opcodes_h_l1259_c2_6935
n8_MUX_uxn_opcodes_h_l1259_c2_6935 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1259_c2_6935_cond,
n8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue,
n8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse,
n8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935
result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935
result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935
result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_cond,
result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935
result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935
result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935
result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935
result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_left,
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_right,
BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output);

-- t8_MUX_uxn_opcodes_h_l1272_c7_61a7
t8_MUX_uxn_opcodes_h_l1272_c7_61a7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond,
t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue,
t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse,
t8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output);

-- n8_MUX_uxn_opcodes_h_l1272_c7_61a7
n8_MUX_uxn_opcodes_h_l1272_c7_61a7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond,
n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue,
n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse,
n8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7
result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_cond,
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149
BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_left,
BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_right,
BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output);

-- t8_MUX_uxn_opcodes_h_l1275_c7_bbc3
t8_MUX_uxn_opcodes_h_l1275_c7_bbc3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond,
t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue,
t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse,
t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output);

-- n8_MUX_uxn_opcodes_h_l1275_c7_bbc3
n8_MUX_uxn_opcodes_h_l1275_c7_bbc3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond,
n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue,
n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse,
n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3
result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3
result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3
result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_left,
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_right,
BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output);

-- n8_MUX_uxn_opcodes_h_l1278_c7_5eb1
n8_MUX_uxn_opcodes_h_l1278_c7_5eb1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond,
n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue,
n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse,
n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2
sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_ins,
sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_x,
sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_y,
sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3
BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_left,
BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_right,
BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_return_output);

-- MUX_uxn_opcodes_h_l1283_c21_7ac7
MUX_uxn_opcodes_h_l1283_c21_7ac7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1283_c21_7ac7_cond,
MUX_uxn_opcodes_h_l1283_c21_7ac7_iftrue,
MUX_uxn_opcodes_h_l1283_c21_7ac7_iffalse,
MUX_uxn_opcodes_h_l1283_c21_7ac7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output,
 t8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
 n8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output,
 t8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output,
 n8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output,
 t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output,
 n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output,
 n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output,
 sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_return_output,
 MUX_uxn_opcodes_h_l1283_c21_7ac7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1264_c3_4979 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1269_c3_0c86 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1273_c3_93b8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1282_c3_d7e5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_439c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_4902_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_e741_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_8b79_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1275_l1278_DUPLICATE_181a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1287_l1255_DUPLICATE_b40d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1273_c3_93b8 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1273_c3_93b8;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1264_c3_4979 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1264_c3_4979;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1269_c3_0c86 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1269_c3_0c86;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1282_c3_d7e5 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1282_c3_d7e5;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse := t8;
     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1259_c2_6935_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1259_c6_8358] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_left;
     BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output := BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1259_c2_6935_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1275_l1278_DUPLICATE_181a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1275_l1278_DUPLICATE_181a_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1283_c21_69e3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1259_c2_6935_return_output := result.is_pc_updated;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_4902 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_4902_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_8b79 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_8b79_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1272_c11_5503] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_left;
     BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output := BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1280_c30_f0f2] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_ins;
     sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_x;
     sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_return_output := sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1275_c11_1149] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_left;
     BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output := BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_e741 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_e741_return_output := result.is_stack_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1259_c2_6935_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_439c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_439c_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1278_c11_f038] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_left;
     BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output := BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1259_c6_8358_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1272_c11_5503_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1275_c11_1149_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1278_c11_f038_return_output;
     VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1283_c21_69e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_4902_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_4902_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_4902_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_8b79_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_8b79_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_8b79_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_e741_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_e741_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1275_l1278_l1272_DUPLICATE_e741_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1275_l1278_DUPLICATE_181a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1275_l1278_DUPLICATE_181a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_439c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_439c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_439c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1275_l1259_l1278_l1272_DUPLICATE_439c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1259_c2_6935_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1259_c2_6935_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1259_c2_6935_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1259_c2_6935_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1280_c30_f0f2_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1278_c7_5eb1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;

     -- t8_MUX[uxn_opcodes_h_l1275_c7_bbc3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond <= VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond;
     t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue;
     t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output := t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1278_c7_5eb1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1278_c7_5eb1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;

     -- MUX[uxn_opcodes_h_l1283_c21_7ac7] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1283_c21_7ac7_cond <= VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_cond;
     MUX_uxn_opcodes_h_l1283_c21_7ac7_iftrue <= VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_iftrue;
     MUX_uxn_opcodes_h_l1283_c21_7ac7_iffalse <= VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_return_output := MUX_uxn_opcodes_h_l1283_c21_7ac7_return_output;

     -- n8_MUX[uxn_opcodes_h_l1278_c7_5eb1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond <= VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond;
     n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue;
     n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output := n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1278_c7_5eb1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue := VAR_MUX_uxn_opcodes_h_l1283_c21_7ac7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;
     -- n8_MUX[uxn_opcodes_h_l1275_c7_bbc3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond <= VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond;
     n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue;
     n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output := n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1278_c7_5eb1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1275_c7_bbc3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1275_c7_bbc3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;

     -- t8_MUX[uxn_opcodes_h_l1272_c7_61a7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond <= VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond;
     t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue;
     t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output := t8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1275_c7_bbc3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1275_c7_bbc3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1278_c7_5eb1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1272_c7_61a7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1275_c7_bbc3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;

     -- t8_MUX[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1259_c2_6935_cond <= VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_cond;
     t8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue;
     t8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output := t8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;

     -- n8_MUX[uxn_opcodes_h_l1272_c7_61a7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond <= VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_cond;
     n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue;
     n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output := n8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1272_c7_61a7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1272_c7_61a7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1272_c7_61a7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1275_c7_bbc3_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1272_c7_61a7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output := result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;

     -- n8_MUX[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1259_c2_6935_cond <= VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_cond;
     n8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue;
     n8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output := n8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1272_c7_61a7_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1259_c2_6935] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_return_output := result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1287_l1255_DUPLICATE_b40d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1287_l1255_DUPLICATE_b40d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_188e(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1259_c2_6935_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1259_c2_6935_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1287_l1255_DUPLICATE_b40d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1287_l1255_DUPLICATE_b40d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
