-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity eor_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_fedec265;
architecture arch of eor_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1136_c6_6d53]
signal BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1136_c2_b196]
signal n8_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1136_c2_b196]
signal t8_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1136_c2_b196]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1136_c2_b196]
signal result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1136_c2_b196]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1136_c2_b196]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1136_c2_b196]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1136_c2_b196]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1141_c11_7eae]
signal BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1141_c7_4f27]
signal n8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1141_c7_4f27]
signal t8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1141_c7_4f27]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1141_c7_4f27]
signal result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1141_c7_4f27]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1141_c7_4f27]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1141_c7_4f27]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1141_c7_4f27]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1144_c11_b81f]
signal BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1144_c7_5bf0]
signal n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1144_c7_5bf0]
signal t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1144_c7_5bf0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1144_c7_5bf0]
signal result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1144_c7_5bf0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1144_c7_5bf0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1144_c7_5bf0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1144_c7_5bf0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1148_c11_ba3d]
signal BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1148_c7_a513]
signal n8_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1148_c7_a513]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1148_c7_a513]
signal result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1148_c7_a513]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1148_c7_a513]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1148_c7_a513]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1148_c7_a513]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1151_c11_4de8]
signal BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1151_c7_e305]
signal n8_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1151_c7_e305]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1151_c7_e305]
signal result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1151_c7_e305]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1151_c7_e305]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1151_c7_e305]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1151_c7_e305]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1154_c30_8cdb]
signal sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1157_c21_d64b]
signal BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1159_c11_2a12]
signal BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1159_c7_78cc]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1159_c7_78cc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1159_c7_78cc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53
BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_left,
BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_right,
BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output);

-- n8_MUX_uxn_opcodes_h_l1136_c2_b196
n8_MUX_uxn_opcodes_h_l1136_c2_b196 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1136_c2_b196_cond,
n8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue,
n8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse,
n8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output);

-- t8_MUX_uxn_opcodes_h_l1136_c2_b196
t8_MUX_uxn_opcodes_h_l1136_c2_b196 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1136_c2_b196_cond,
t8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue,
t8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse,
t8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196
result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_cond,
result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196
result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196
result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196
result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196
result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae
BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_left,
BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_right,
BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output);

-- n8_MUX_uxn_opcodes_h_l1141_c7_4f27
n8_MUX_uxn_opcodes_h_l1141_c7_4f27 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond,
n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue,
n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse,
n8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output);

-- t8_MUX_uxn_opcodes_h_l1141_c7_4f27
t8_MUX_uxn_opcodes_h_l1141_c7_4f27 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond,
t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue,
t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse,
t8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27
result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_cond,
result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27
result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27
result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27
result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27
result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f
BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_left,
BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_right,
BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output);

-- n8_MUX_uxn_opcodes_h_l1144_c7_5bf0
n8_MUX_uxn_opcodes_h_l1144_c7_5bf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond,
n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue,
n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse,
n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output);

-- t8_MUX_uxn_opcodes_h_l1144_c7_5bf0
t8_MUX_uxn_opcodes_h_l1144_c7_5bf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond,
t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue,
t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse,
t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0
result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0
result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0
result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0
result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d
BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_left,
BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_right,
BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output);

-- n8_MUX_uxn_opcodes_h_l1148_c7_a513
n8_MUX_uxn_opcodes_h_l1148_c7_a513 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1148_c7_a513_cond,
n8_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue,
n8_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse,
n8_MUX_uxn_opcodes_h_l1148_c7_a513_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513
result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_cond,
result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513
result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513
result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513
result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513
result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8
BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_left,
BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_right,
BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output);

-- n8_MUX_uxn_opcodes_h_l1151_c7_e305
n8_MUX_uxn_opcodes_h_l1151_c7_e305 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1151_c7_e305_cond,
n8_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue,
n8_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse,
n8_MUX_uxn_opcodes_h_l1151_c7_e305_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305
result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_cond,
result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305
result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305
result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305
result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305
result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb
sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_ins,
sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_x,
sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_y,
sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b
BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_left,
BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_right,
BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12
BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_left,
BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_right,
BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc
result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc
result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc
result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output,
 n8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
 t8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output,
 n8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output,
 t8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output,
 n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output,
 t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output,
 n8_MUX_uxn_opcodes_h_l1148_c7_a513_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output,
 n8_MUX_uxn_opcodes_h_l1151_c7_e305_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output,
 sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1138_c3_9ef8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1142_c3_3830 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1146_c3_c766 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1149_c3_3a7f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1156_c3_31b0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1151_c7_e305_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_37d0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_641e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_a080_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_8135_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1159_DUPLICATE_add5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1132_l1165_DUPLICATE_257d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1156_c3_31b0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1156_c3_31b0;
     VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1146_c3_c766 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1146_c3_c766;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1142_c3_3830 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1142_c3_3830;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1149_c3_3a7f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1149_c3_3a7f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1138_c3_9ef8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1138_c3_9ef8;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l1154_c30_8cdb] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_ins;
     sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_x;
     sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_return_output := sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1148_c11_ba3d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1151_c11_4de8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_a080 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_a080_return_output := result.sp_relative_shift;

     -- BIN_OP_XOR[uxn_opcodes_h_l1157_c21_d64b] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_left;
     BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_return_output := BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1151_c7_e305] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1151_c7_e305_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1136_c6_6d53] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_left;
     BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output := BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1159_c11_2a12] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_left;
     BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_return_output := BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1141_c11_7eae] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_left;
     BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output := BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1144_c11_b81f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_641e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_641e_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_8135 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_8135_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_37d0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_37d0_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1159_DUPLICATE_add5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1159_DUPLICATE_add5_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1136_c6_6d53_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1141_c11_7eae_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1144_c11_b81f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1148_c11_ba3d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1151_c11_4de8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c11_2a12_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1157_c21_d64b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_a080_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_a080_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_a080_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_a080_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_a080_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1159_DUPLICATE_add5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1159_DUPLICATE_add5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1159_DUPLICATE_add5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1159_DUPLICATE_add5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1159_DUPLICATE_add5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_8135_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_8135_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_8135_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_8135_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_8135_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_641e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_641e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_641e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_641e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1148_l1144_l1141_l1136_l1159_DUPLICATE_641e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_37d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_37d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_37d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_37d0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1151_l1148_l1144_l1141_l1136_DUPLICATE_37d0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1151_c7_e305_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1154_c30_8cdb_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1151_c7_e305] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;

     -- t8_MUX[uxn_opcodes_h_l1144_c7_5bf0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond <= VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond;
     t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue;
     t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output := t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1159_c7_78cc] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1151_c7_e305] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_return_output := result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1159_c7_78cc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1159_c7_78cc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1151_c7_e305] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;

     -- n8_MUX[uxn_opcodes_h_l1151_c7_e305] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1151_c7_e305_cond <= VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_cond;
     n8_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue;
     n8_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_return_output := n8_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1159_c7_78cc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1151_c7_e305] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1148_c7_a513] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1151_c7_e305] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;

     -- t8_MUX[uxn_opcodes_h_l1141_c7_4f27] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond <= VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond;
     t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue;
     t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output := t8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1151_c7_e305] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;

     -- n8_MUX[uxn_opcodes_h_l1148_c7_a513] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1148_c7_a513_cond <= VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_cond;
     n8_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue;
     n8_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_return_output := n8_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1148_c7_a513] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1148_c7_a513] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_return_output := result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1151_c7_e305_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;
     -- n8_MUX[uxn_opcodes_h_l1144_c7_5bf0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond <= VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond;
     n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue;
     n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output := n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1144_c7_5bf0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1148_c7_a513] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1144_c7_5bf0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1148_c7_a513] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1148_c7_a513] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1144_c7_5bf0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;

     -- t8_MUX[uxn_opcodes_h_l1136_c2_b196] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1136_c2_b196_cond <= VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_cond;
     t8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue;
     t8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output := t8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1148_c7_a513_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1144_c7_5bf0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1141_c7_4f27] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output := result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1144_c7_5bf0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;

     -- n8_MUX[uxn_opcodes_h_l1141_c7_4f27] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond <= VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_cond;
     n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue;
     n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output := n8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1141_c7_4f27] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1141_c7_4f27] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1144_c7_5bf0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1144_c7_5bf0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1136_c2_b196] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1136_c2_b196] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1141_c7_4f27] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;

     -- n8_MUX[uxn_opcodes_h_l1136_c2_b196] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1136_c2_b196_cond <= VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_cond;
     n8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue;
     n8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output := n8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1141_c7_4f27] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1136_c2_b196] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_return_output := result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1141_c7_4f27] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1136_c2_b196_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1141_c7_4f27_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1136_c2_b196] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1136_c2_b196] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1136_c2_b196] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1132_l1165_DUPLICATE_257d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1132_l1165_DUPLICATE_257d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1136_c2_b196_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1132_l1165_DUPLICATE_257d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1132_l1165_DUPLICATE_257d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
